magic
tech sky130A
magscale 1 2
timestamp 1647860640
<< viali >>
rect 2237 11305 2271 11339
rect 4169 11305 4203 11339
rect 5273 11305 5307 11339
rect 5917 11305 5951 11339
rect 6469 11305 6503 11339
rect 9229 11305 9263 11339
rect 1777 11237 1811 11271
rect 3433 11237 3467 11271
rect 4537 11237 4571 11271
rect 7665 11237 7699 11271
rect 9137 11237 9171 11271
rect 9505 11237 9539 11271
rect 4629 11169 4663 11203
rect 5825 11169 5859 11203
rect 6653 11169 6687 11203
rect 8769 11169 8803 11203
rect 2053 11101 2087 11135
rect 2421 11101 2455 11135
rect 2605 11101 2639 11135
rect 2789 11101 2823 11135
rect 3617 11101 3651 11135
rect 3893 11101 3927 11135
rect 4353 11101 4387 11135
rect 5089 11101 5123 11135
rect 6193 11101 6227 11135
rect 6837 11101 6871 11135
rect 7205 11101 7239 11135
rect 7481 11101 7515 11135
rect 2881 11033 2915 11067
rect 3065 11033 3099 11067
rect 3249 11033 3283 11067
rect 3985 11033 4019 11067
rect 5457 11033 5491 11067
rect 5641 11033 5675 11067
rect 6377 11033 6411 11067
rect 6929 11033 6963 11067
rect 7297 11033 7331 11067
rect 7757 11033 7791 11067
rect 8033 11033 8067 11067
rect 8217 11033 8251 11067
rect 1961 10965 1995 10999
rect 3801 10965 3835 10999
rect 4905 10965 4939 10999
rect 8401 10965 8435 10999
rect 8493 10965 8527 10999
rect 4445 10761 4479 10795
rect 5089 10761 5123 10795
rect 5641 10761 5675 10795
rect 7849 10761 7883 10795
rect 1685 10693 1719 10727
rect 1501 10625 1535 10659
rect 1777 10625 1811 10659
rect 3617 10625 3651 10659
rect 4905 10625 4939 10659
rect 5181 10625 5215 10659
rect 6009 10625 6043 10659
rect 6193 10625 6227 10659
rect 6929 10625 6963 10659
rect 7113 10625 7147 10659
rect 7205 10625 7239 10659
rect 7665 10625 7699 10659
rect 7941 10625 7975 10659
rect 8309 10625 8343 10659
rect 9321 10625 9355 10659
rect 1317 10557 1351 10591
rect 2145 10557 2179 10591
rect 4181 10557 4215 10591
rect 9413 10557 9447 10591
rect 6653 10489 6687 10523
rect 8493 10489 8527 10523
rect 4813 10421 4847 10455
rect 5273 10421 5307 10455
rect 5825 10421 5859 10455
rect 6285 10421 6319 10455
rect 7297 10421 7331 10455
rect 7481 10421 7515 10455
rect 8125 10421 8159 10455
rect 8677 10421 8711 10455
rect 4445 10217 4479 10251
rect 8769 10217 8803 10251
rect 2697 10149 2731 10183
rect 3617 10149 3651 10183
rect 8493 10149 8527 10183
rect 1317 10081 1351 10115
rect 8309 10081 8343 10115
rect 1961 10013 1995 10047
rect 2053 10013 2087 10047
rect 3433 10013 3467 10047
rect 3801 10013 3835 10047
rect 5733 10013 5767 10047
rect 6469 10013 6503 10047
rect 7941 10013 7975 10047
rect 8585 10013 8619 10047
rect 9413 10013 9447 10047
rect 2789 9945 2823 9979
rect 5909 9877 5943 9911
rect 9505 9673 9539 9707
rect 1501 9605 1535 9639
rect 3341 9537 3375 9571
rect 3433 9537 3467 9571
rect 5273 9537 5307 9571
rect 6377 9537 6411 9571
rect 6561 9537 6595 9571
rect 6837 9537 6871 9571
rect 8677 9537 8711 9571
rect 1225 9469 1259 9503
rect 3801 9469 3835 9503
rect 7205 9469 7239 9503
rect 6193 9401 6227 9435
rect 6745 9401 6779 9435
rect 2973 9333 3007 9367
rect 3157 9333 3191 9367
rect 5837 9333 5871 9367
rect 9237 9333 9271 9367
rect 1685 9129 1719 9163
rect 2329 9129 2363 9163
rect 2789 9129 2823 9163
rect 3157 9129 3191 9163
rect 3985 9129 4019 9163
rect 9413 9129 9447 9163
rect 4905 9061 4939 9095
rect 5273 9061 5307 9095
rect 5733 9061 5767 9095
rect 6101 9061 6135 9095
rect 2513 8993 2547 9027
rect 8033 8993 8067 9027
rect 1501 8925 1535 8959
rect 1961 8925 1995 8959
rect 2053 8925 2087 8959
rect 2697 8925 2731 8959
rect 3617 8925 3651 8959
rect 4261 8925 4295 8959
rect 4537 8925 4571 8959
rect 5181 8925 5215 8959
rect 5457 8925 5491 8959
rect 5549 8925 5583 8959
rect 5917 8925 5951 8959
rect 8309 8925 8343 8959
rect 8769 8925 8803 8959
rect 1317 8857 1351 8891
rect 3433 8857 3467 8891
rect 4077 8857 4111 8891
rect 4721 8857 4755 8891
rect 7757 8857 7791 8891
rect 1869 8789 1903 8823
rect 3801 8789 3835 8823
rect 4445 8789 4479 8823
rect 4997 8789 5031 8823
rect 6285 8789 6319 8823
rect 8217 8789 8251 8823
rect 8493 8789 8527 8823
rect 1593 8585 1627 8619
rect 6009 8585 6043 8619
rect 7205 8585 7239 8619
rect 9413 8585 9447 8619
rect 5457 8517 5491 8551
rect 5641 8517 5675 8551
rect 5825 8517 5859 8551
rect 1685 8449 1719 8483
rect 1777 8449 1811 8483
rect 3617 8449 3651 8483
rect 4353 8449 4387 8483
rect 4997 8449 5031 8483
rect 5181 8449 5215 8483
rect 6285 8449 6319 8483
rect 6561 8449 6595 8483
rect 9137 8449 9171 8483
rect 9229 8449 9263 8483
rect 1409 8381 1443 8415
rect 2145 8381 2179 8415
rect 4813 8381 4847 8415
rect 7389 8381 7423 8415
rect 8861 8381 8895 8415
rect 5365 8313 5399 8347
rect 4181 8245 4215 8279
rect 4629 8245 4663 8279
rect 6377 8245 6411 8279
rect 2697 8041 2731 8075
rect 6009 8041 6043 8075
rect 9413 8041 9447 8075
rect 5733 7973 5767 8007
rect 6101 7905 6135 7939
rect 1961 7837 1995 7871
rect 2053 7837 2087 7871
rect 2789 7837 2823 7871
rect 4261 7837 4295 7871
rect 4353 7837 4387 7871
rect 5089 7837 5123 7871
rect 5825 7837 5859 7871
rect 8217 7837 8251 7871
rect 8585 7837 8619 7871
rect 8769 7837 8803 7871
rect 1317 7769 1351 7803
rect 3433 7769 3467 7803
rect 3617 7769 3651 7803
rect 6377 7769 6411 7803
rect 4997 7701 5031 7735
rect 7849 7701 7883 7735
rect 8125 7701 8159 7735
rect 8309 7701 8343 7735
rect 8401 7701 8435 7735
rect 1317 7497 1351 7531
rect 1409 7497 1443 7531
rect 5929 7497 5963 7531
rect 3525 7361 3559 7395
rect 3893 7361 3927 7395
rect 5365 7361 5399 7395
rect 6377 7361 6411 7395
rect 8217 7361 8251 7395
rect 8953 7361 8987 7395
rect 3157 7293 3191 7327
rect 3433 7293 3467 7327
rect 6745 7293 6779 7327
rect 6193 7225 6227 7259
rect 1685 7157 1719 7191
rect 8401 7157 8435 7191
rect 8781 7157 8815 7191
rect 9045 7157 9079 7191
rect 9413 7157 9447 7191
rect 2807 6953 2841 6987
rect 5733 6885 5767 6919
rect 3065 6817 3099 6851
rect 6285 6817 6319 6851
rect 3249 6749 3283 6783
rect 4261 6749 4295 6783
rect 4353 6749 4387 6783
rect 5089 6749 5123 6783
rect 6009 6749 6043 6783
rect 7849 6749 7883 6783
rect 8585 6749 8619 6783
rect 9505 6749 9539 6783
rect 3617 6681 3651 6715
rect 8861 6681 8895 6715
rect 1317 6613 1351 6647
rect 3433 6613 3467 6647
rect 4997 6613 5031 6647
rect 5825 6613 5859 6647
rect 7941 6613 7975 6647
rect 5917 6409 5951 6443
rect 1593 6341 1627 6375
rect 7665 6341 7699 6375
rect 3249 6273 3283 6307
rect 5089 6273 5123 6307
rect 6009 6273 6043 6307
rect 6377 6273 6411 6307
rect 6561 6273 6595 6307
rect 6745 6273 6779 6307
rect 7021 6273 7055 6307
rect 7297 6273 7331 6307
rect 7389 6273 7423 6307
rect 9505 6273 9539 6307
rect 1317 6205 1351 6239
rect 3617 6205 3651 6239
rect 6929 6205 6963 6239
rect 6193 6137 6227 6171
rect 9321 6137 9355 6171
rect 3065 6069 3099 6103
rect 5653 6069 5687 6103
rect 9137 6069 9171 6103
rect 3709 5865 3743 5899
rect 4077 5865 4111 5899
rect 5549 5865 5583 5899
rect 6285 5865 6319 5899
rect 6929 5865 6963 5899
rect 7757 5865 7791 5899
rect 8861 5865 8895 5899
rect 6653 5797 6687 5831
rect 1593 5729 1627 5763
rect 7297 5729 7331 5763
rect 9229 5729 9263 5763
rect 1317 5661 1351 5695
rect 4169 5661 4203 5695
rect 4261 5661 4295 5695
rect 6193 5661 6227 5695
rect 6837 5661 6871 5695
rect 7481 5661 7515 5695
rect 7757 5661 7791 5695
rect 8125 5661 8159 5695
rect 8309 5661 8343 5695
rect 8585 5661 8619 5695
rect 9045 5661 9079 5695
rect 9321 5661 9355 5695
rect 1869 5593 1903 5627
rect 1501 5525 1535 5559
rect 3341 5525 3375 5559
rect 7665 5525 7699 5559
rect 9413 5525 9447 5559
rect 4813 5321 4847 5355
rect 5733 5321 5767 5355
rect 9321 5321 9355 5355
rect 5089 5253 5123 5287
rect 7021 5253 7055 5287
rect 7757 5253 7791 5287
rect 8493 5253 8527 5287
rect 8861 5253 8895 5287
rect 3433 5185 3467 5219
rect 4077 5185 4111 5219
rect 4169 5185 4203 5219
rect 7113 5185 7147 5219
rect 7941 5185 7975 5219
rect 8309 5185 8343 5219
rect 8953 5185 8987 5219
rect 9229 5185 9263 5219
rect 9505 5185 9539 5219
rect 8125 5117 8159 5151
rect 4905 5049 4939 5083
rect 8677 5049 8711 5083
rect 7205 4981 7239 5015
rect 7573 4981 7607 5015
rect 3433 4777 3467 4811
rect 4445 4777 4479 4811
rect 5089 4777 5123 4811
rect 5825 4777 5859 4811
rect 9137 4777 9171 4811
rect 5549 4709 5583 4743
rect 6837 4641 6871 4675
rect 4077 4573 4111 4607
rect 4721 4573 4755 4607
rect 5365 4573 5399 4607
rect 5733 4573 5767 4607
rect 6469 4573 6503 4607
rect 8309 4573 8343 4607
rect 9321 4573 9355 4607
rect 9413 4573 9447 4607
rect 8873 4505 8907 4539
rect 4261 4437 4295 4471
rect 4905 4437 4939 4471
rect 6193 4437 6227 4471
rect 3341 4233 3375 4267
rect 8769 4233 8803 4267
rect 3801 4165 3835 4199
rect 7113 4165 7147 4199
rect 8493 4165 8527 4199
rect 9137 4165 9171 4199
rect 3525 4097 3559 4131
rect 3985 4097 4019 4131
rect 4169 4097 4203 4131
rect 6285 4097 6319 4131
rect 7389 4097 7423 4131
rect 7665 4097 7699 4131
rect 8125 4097 8159 4131
rect 8677 4097 8711 4131
rect 8953 4097 8987 4131
rect 9505 4097 9539 4131
rect 4445 4029 4479 4063
rect 4813 4029 4847 4063
rect 7481 4029 7515 4063
rect 8309 4029 8343 4063
rect 7849 3961 7883 3995
rect 9321 3961 9355 3995
rect 3709 3893 3743 3927
rect 4261 3893 4295 3927
rect 6845 3893 6879 3927
rect 7205 3893 7239 3927
rect 7941 3893 7975 3927
rect 3617 3689 3651 3723
rect 5365 3689 5399 3723
rect 6285 3689 6319 3723
rect 8777 3689 8811 3723
rect 9505 3689 9539 3723
rect 4721 3621 4755 3655
rect 3433 3485 3467 3519
rect 3709 3485 3743 3519
rect 3985 3485 4019 3519
rect 4261 3485 4295 3519
rect 4537 3485 4571 3519
rect 4997 3485 5031 3519
rect 5733 3485 5767 3519
rect 6377 3485 6411 3519
rect 6745 3485 6779 3519
rect 8217 3485 8251 3519
rect 9137 3485 9171 3519
rect 5089 3417 5123 3451
rect 5273 3417 5307 3451
rect 5917 3417 5951 3451
rect 6101 3417 6135 3451
rect 9229 3417 9263 3451
rect 3893 3349 3927 3383
rect 4169 3349 4203 3383
rect 4445 3349 4479 3383
rect 4905 3349 4939 3383
rect 8953 3349 8987 3383
rect 8033 3145 8067 3179
rect 8309 3145 8343 3179
rect 6561 3077 6595 3111
rect 3433 3009 3467 3043
rect 3709 3009 3743 3043
rect 5549 3009 5583 3043
rect 6285 3009 6319 3043
rect 8953 3009 8987 3043
rect 9045 3009 9079 3043
rect 9505 3009 9539 3043
rect 4077 2941 4111 2975
rect 3617 2873 3651 2907
rect 9413 2873 9447 2907
rect 6113 2805 6147 2839
rect 9229 2805 9263 2839
rect 5917 2601 5951 2635
rect 8409 2601 8443 2635
rect 5457 2465 5491 2499
rect 6009 2465 6043 2499
rect 9045 2465 9079 2499
rect 3341 2397 3375 2431
rect 5365 2397 5399 2431
rect 5733 2397 5767 2431
rect 6377 2397 6411 2431
rect 7849 2397 7883 2431
rect 3617 2329 3651 2363
rect 9229 2329 9263 2363
rect 9321 2329 9355 2363
rect 5089 2261 5123 2295
rect 8309 2057 8343 2091
rect 8585 2057 8619 2091
rect 9045 2057 9079 2091
rect 3525 1989 3559 2023
rect 3709 1989 3743 2023
rect 3893 1989 3927 2023
rect 4353 1989 4387 2023
rect 4629 1921 4663 1955
rect 6561 1921 6595 1955
rect 8125 1921 8159 1955
rect 8861 1921 8895 1955
rect 8953 1921 8987 1955
rect 4905 1853 4939 1887
rect 6377 1853 6411 1887
rect 9413 1853 9447 1887
rect 8033 1785 8067 1819
rect 4077 1717 4111 1751
rect 4445 1717 4479 1751
rect 9229 1717 9263 1751
rect 5089 1513 5123 1547
rect 6469 1513 6503 1547
rect 8033 1513 8067 1547
rect 9229 1513 9263 1547
rect 5549 1445 5583 1479
rect 3341 1377 3375 1411
rect 3617 1377 3651 1411
rect 5365 1309 5399 1343
rect 5733 1309 5767 1343
rect 7113 1309 7147 1343
rect 7205 1309 7239 1343
rect 6377 1241 6411 1275
rect 7849 1241 7883 1275
rect 8309 1173 8343 1207
rect 8493 1173 8527 1207
rect 8677 1173 8711 1207
rect 8861 1173 8895 1207
rect 9321 1173 9355 1207
<< metal1 >>
rect 2774 11568 2780 11620
rect 2832 11608 2838 11620
rect 4246 11608 4252 11620
rect 2832 11580 4252 11608
rect 2832 11568 2838 11580
rect 4246 11568 4252 11580
rect 4304 11568 4310 11620
rect 1854 11500 1860 11552
rect 1912 11540 1918 11552
rect 4982 11540 4988 11552
rect 1912 11512 4988 11540
rect 1912 11500 1918 11512
rect 4982 11500 4988 11512
rect 5040 11500 5046 11552
rect 920 11450 9844 11472
rect 920 11398 2566 11450
rect 2618 11398 2630 11450
rect 2682 11398 2694 11450
rect 2746 11398 2758 11450
rect 2810 11398 2822 11450
rect 2874 11398 7566 11450
rect 7618 11398 7630 11450
rect 7682 11398 7694 11450
rect 7746 11398 7758 11450
rect 7810 11398 7822 11450
rect 7874 11398 9844 11450
rect 920 11376 9844 11398
rect 1394 11296 1400 11348
rect 1452 11336 1458 11348
rect 2225 11339 2283 11345
rect 2225 11336 2237 11339
rect 1452 11308 2237 11336
rect 1452 11296 1458 11308
rect 2225 11305 2237 11308
rect 2271 11336 2283 11339
rect 2406 11336 2412 11348
rect 2271 11308 2412 11336
rect 2271 11305 2283 11308
rect 2225 11299 2283 11305
rect 2406 11296 2412 11308
rect 2464 11296 2470 11348
rect 4157 11339 4215 11345
rect 4157 11336 4169 11339
rect 2608 11308 4169 11336
rect 1765 11271 1823 11277
rect 1765 11237 1777 11271
rect 1811 11268 1823 11271
rect 1854 11268 1860 11280
rect 1811 11240 1860 11268
rect 1811 11237 1823 11240
rect 1765 11231 1823 11237
rect 1854 11228 1860 11240
rect 1912 11228 1918 11280
rect 2314 11228 2320 11280
rect 2372 11268 2378 11280
rect 2608 11268 2636 11308
rect 4157 11305 4169 11308
rect 4203 11305 4215 11339
rect 4157 11299 4215 11305
rect 2372 11240 2636 11268
rect 2372 11228 2378 11240
rect 2958 11228 2964 11280
rect 3016 11268 3022 11280
rect 3421 11271 3479 11277
rect 3421 11268 3433 11271
rect 3016 11240 3433 11268
rect 3016 11228 3022 11240
rect 3421 11237 3433 11240
rect 3467 11268 3479 11271
rect 3510 11268 3516 11280
rect 3467 11240 3516 11268
rect 3467 11237 3479 11240
rect 3421 11231 3479 11237
rect 3510 11228 3516 11240
rect 3568 11228 3574 11280
rect 4172 11200 4200 11299
rect 4614 11296 4620 11348
rect 4672 11336 4678 11348
rect 5261 11339 5319 11345
rect 5261 11336 5273 11339
rect 4672 11308 5273 11336
rect 4672 11296 4678 11308
rect 5261 11305 5273 11308
rect 5307 11336 5319 11339
rect 5442 11336 5448 11348
rect 5307 11308 5448 11336
rect 5307 11305 5319 11308
rect 5261 11299 5319 11305
rect 5442 11296 5448 11308
rect 5500 11296 5506 11348
rect 5626 11296 5632 11348
rect 5684 11336 5690 11348
rect 5905 11339 5963 11345
rect 5905 11336 5917 11339
rect 5684 11308 5917 11336
rect 5684 11296 5690 11308
rect 5905 11305 5917 11308
rect 5951 11305 5963 11339
rect 5905 11299 5963 11305
rect 6457 11339 6515 11345
rect 6457 11305 6469 11339
rect 6503 11336 6515 11339
rect 8110 11336 8116 11348
rect 6503 11308 8116 11336
rect 6503 11305 6515 11308
rect 6457 11299 6515 11305
rect 8110 11296 8116 11308
rect 8168 11296 8174 11348
rect 8662 11296 8668 11348
rect 8720 11336 8726 11348
rect 9217 11339 9275 11345
rect 9217 11336 9229 11339
rect 8720 11308 9229 11336
rect 8720 11296 8726 11308
rect 9217 11305 9229 11308
rect 9263 11305 9275 11339
rect 9217 11299 9275 11305
rect 4522 11268 4528 11280
rect 4483 11240 4528 11268
rect 4522 11228 4528 11240
rect 4580 11228 4586 11280
rect 5074 11228 5080 11280
rect 5132 11268 5138 11280
rect 7653 11271 7711 11277
rect 5132 11240 6224 11268
rect 5132 11228 5138 11240
rect 4614 11200 4620 11212
rect 2056 11172 3924 11200
rect 4172 11172 4620 11200
rect 1670 11092 1676 11144
rect 1728 11132 1734 11144
rect 2056 11141 2084 11172
rect 2041 11135 2099 11141
rect 2041 11132 2053 11135
rect 1728 11104 2053 11132
rect 1728 11092 1734 11104
rect 2041 11101 2053 11104
rect 2087 11101 2099 11135
rect 2406 11132 2412 11144
rect 2367 11104 2412 11132
rect 2041 11095 2099 11101
rect 2406 11092 2412 11104
rect 2464 11092 2470 11144
rect 2593 11135 2651 11141
rect 2593 11101 2605 11135
rect 2639 11132 2651 11135
rect 2682 11132 2688 11144
rect 2639 11104 2688 11132
rect 2639 11101 2651 11104
rect 2593 11095 2651 11101
rect 2682 11092 2688 11104
rect 2740 11092 2746 11144
rect 3896 11141 3924 11172
rect 4614 11160 4620 11172
rect 4672 11160 4678 11212
rect 5813 11203 5871 11209
rect 5813 11169 5825 11203
rect 5859 11200 5871 11203
rect 5902 11200 5908 11212
rect 5859 11172 5908 11200
rect 5859 11169 5871 11172
rect 5813 11163 5871 11169
rect 5902 11160 5908 11172
rect 5960 11160 5966 11212
rect 6196 11200 6224 11240
rect 7653 11237 7665 11271
rect 7699 11268 7711 11271
rect 7926 11268 7932 11280
rect 7699 11240 7932 11268
rect 7699 11237 7711 11240
rect 7653 11231 7711 11237
rect 7926 11228 7932 11240
rect 7984 11228 7990 11280
rect 9125 11271 9183 11277
rect 9125 11237 9137 11271
rect 9171 11268 9183 11271
rect 9493 11271 9551 11277
rect 9493 11268 9505 11271
rect 9171 11240 9505 11268
rect 9171 11237 9183 11240
rect 9125 11231 9183 11237
rect 9493 11237 9505 11240
rect 9539 11268 9551 11271
rect 16574 11268 16580 11280
rect 9539 11240 16580 11268
rect 9539 11237 9551 11240
rect 9493 11231 9551 11237
rect 16574 11228 16580 11240
rect 16632 11228 16638 11280
rect 6641 11203 6699 11209
rect 6641 11200 6653 11203
rect 6196 11172 6653 11200
rect 6196 11144 6224 11172
rect 6641 11169 6653 11172
rect 6687 11169 6699 11203
rect 6641 11163 6699 11169
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 8757 11203 8815 11209
rect 8757 11200 8769 11203
rect 7156 11172 8769 11200
rect 7156 11160 7162 11172
rect 8757 11169 8769 11172
rect 8803 11169 8815 11203
rect 8757 11163 8815 11169
rect 2777 11135 2835 11141
rect 2777 11101 2789 11135
rect 2823 11132 2835 11135
rect 3605 11135 3663 11141
rect 3605 11132 3617 11135
rect 2823 11104 3617 11132
rect 2823 11101 2835 11104
rect 2777 11095 2835 11101
rect 3605 11101 3617 11104
rect 3651 11101 3663 11135
rect 3605 11095 3663 11101
rect 3881 11135 3939 11141
rect 3881 11101 3893 11135
rect 3927 11101 3939 11135
rect 4338 11132 4344 11144
rect 4299 11104 4344 11132
rect 3881 11095 3939 11101
rect 4338 11092 4344 11104
rect 4396 11092 4402 11144
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11132 5135 11135
rect 6086 11132 6092 11144
rect 5123 11104 6092 11132
rect 5123 11101 5135 11104
rect 5077 11095 5135 11101
rect 6086 11092 6092 11104
rect 6144 11092 6150 11144
rect 6178 11092 6184 11144
rect 6236 11132 6242 11144
rect 6236 11104 6329 11132
rect 6236 11092 6242 11104
rect 6454 11092 6460 11144
rect 6512 11132 6518 11144
rect 6825 11135 6883 11141
rect 6825 11132 6837 11135
rect 6512 11104 6837 11132
rect 6512 11092 6518 11104
rect 6825 11101 6837 11104
rect 6871 11101 6883 11135
rect 7190 11132 7196 11144
rect 7151 11104 7196 11132
rect 6825 11095 6883 11101
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7469 11135 7527 11141
rect 7469 11101 7481 11135
rect 7515 11132 7527 11135
rect 7558 11132 7564 11144
rect 7515 11104 7564 11132
rect 7515 11101 7527 11104
rect 7469 11095 7527 11101
rect 7558 11092 7564 11104
rect 7616 11092 7622 11144
rect 2869 11067 2927 11073
rect 2869 11064 2881 11067
rect 2700 11036 2881 11064
rect 1946 10996 1952 11008
rect 1907 10968 1952 10996
rect 1946 10956 1952 10968
rect 2004 10956 2010 11008
rect 2130 10956 2136 11008
rect 2188 10996 2194 11008
rect 2700 10996 2728 11036
rect 2869 11033 2881 11036
rect 2915 11064 2927 11067
rect 2958 11064 2964 11076
rect 2915 11036 2964 11064
rect 2915 11033 2927 11036
rect 2869 11027 2927 11033
rect 2958 11024 2964 11036
rect 3016 11024 3022 11076
rect 3050 11024 3056 11076
rect 3108 11064 3114 11076
rect 3234 11064 3240 11076
rect 3108 11036 3153 11064
rect 3195 11036 3240 11064
rect 3108 11024 3114 11036
rect 3234 11024 3240 11036
rect 3292 11024 3298 11076
rect 3418 11024 3424 11076
rect 3476 11064 3482 11076
rect 3973 11067 4031 11073
rect 3973 11064 3985 11067
rect 3476 11036 3985 11064
rect 3476 11024 3482 11036
rect 3973 11033 3985 11036
rect 4019 11033 4031 11067
rect 5442 11064 5448 11076
rect 5403 11036 5448 11064
rect 3973 11027 4031 11033
rect 5442 11024 5448 11036
rect 5500 11024 5506 11076
rect 5629 11067 5687 11073
rect 5629 11033 5641 11067
rect 5675 11064 5687 11067
rect 5718 11064 5724 11076
rect 5675 11036 5724 11064
rect 5675 11033 5687 11036
rect 5629 11027 5687 11033
rect 5718 11024 5724 11036
rect 5776 11064 5782 11076
rect 6365 11067 6423 11073
rect 6365 11064 6377 11067
rect 5776 11036 6377 11064
rect 5776 11024 5782 11036
rect 6365 11033 6377 11036
rect 6411 11033 6423 11067
rect 6914 11064 6920 11076
rect 6875 11036 6920 11064
rect 6365 11027 6423 11033
rect 6914 11024 6920 11036
rect 6972 11024 6978 11076
rect 7006 11024 7012 11076
rect 7064 11064 7070 11076
rect 7285 11067 7343 11073
rect 7285 11064 7297 11067
rect 7064 11036 7297 11064
rect 7064 11024 7070 11036
rect 7285 11033 7297 11036
rect 7331 11033 7343 11067
rect 7285 11027 7343 11033
rect 7374 11024 7380 11076
rect 7432 11064 7438 11076
rect 7745 11067 7803 11073
rect 7745 11064 7757 11067
rect 7432 11036 7757 11064
rect 7432 11024 7438 11036
rect 7745 11033 7757 11036
rect 7791 11033 7803 11067
rect 8018 11064 8024 11076
rect 7979 11036 8024 11064
rect 7745 11027 7803 11033
rect 8018 11024 8024 11036
rect 8076 11024 8082 11076
rect 8205 11067 8263 11073
rect 8205 11033 8217 11067
rect 8251 11064 8263 11067
rect 8251 11036 8432 11064
rect 8251 11033 8263 11036
rect 8205 11027 8263 11033
rect 8404 11008 8432 11036
rect 2188 10968 2728 10996
rect 2188 10956 2194 10968
rect 3602 10956 3608 11008
rect 3660 10996 3666 11008
rect 3789 10999 3847 11005
rect 3789 10996 3801 10999
rect 3660 10968 3801 10996
rect 3660 10956 3666 10968
rect 3789 10965 3801 10968
rect 3835 10965 3847 10999
rect 4890 10996 4896 11008
rect 4851 10968 4896 10996
rect 3789 10959 3847 10965
rect 4890 10956 4896 10968
rect 4948 10956 4954 11008
rect 6178 10956 6184 11008
rect 6236 10996 6242 11008
rect 7834 10996 7840 11008
rect 6236 10968 7840 10996
rect 6236 10956 6242 10968
rect 7834 10956 7840 10968
rect 7892 10956 7898 11008
rect 8386 10996 8392 11008
rect 8347 10968 8392 10996
rect 8386 10956 8392 10968
rect 8444 10996 8450 11008
rect 8481 10999 8539 11005
rect 8481 10996 8493 10999
rect 8444 10968 8493 10996
rect 8444 10956 8450 10968
rect 8481 10965 8493 10968
rect 8527 10965 8539 10999
rect 8481 10959 8539 10965
rect 920 10906 9844 10928
rect 920 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 5194 10906
rect 5246 10854 5258 10906
rect 5310 10854 5322 10906
rect 5374 10854 9844 10906
rect 920 10832 9844 10854
rect 4338 10752 4344 10804
rect 4396 10792 4402 10804
rect 4433 10795 4491 10801
rect 4433 10792 4445 10795
rect 4396 10764 4445 10792
rect 4396 10752 4402 10764
rect 4433 10761 4445 10764
rect 4479 10761 4491 10795
rect 4433 10755 4491 10761
rect 5077 10795 5135 10801
rect 5077 10761 5089 10795
rect 5123 10792 5135 10795
rect 5442 10792 5448 10804
rect 5123 10764 5448 10792
rect 5123 10761 5135 10764
rect 5077 10755 5135 10761
rect 3240 10736 3292 10742
rect 1670 10724 1676 10736
rect 1631 10696 1676 10724
rect 1670 10684 1676 10696
rect 1728 10684 1734 10736
rect 3240 10678 3292 10684
rect 1486 10656 1492 10668
rect 1447 10628 1492 10656
rect 1486 10616 1492 10628
rect 1544 10616 1550 10668
rect 1765 10659 1823 10665
rect 1765 10625 1777 10659
rect 1811 10656 1823 10659
rect 1946 10656 1952 10668
rect 1811 10628 1952 10656
rect 1811 10625 1823 10628
rect 1765 10619 1823 10625
rect 1946 10616 1952 10628
rect 2004 10616 2010 10668
rect 3602 10656 3608 10668
rect 3563 10628 3608 10656
rect 3602 10616 3608 10628
rect 3660 10616 3666 10668
rect 4614 10616 4620 10668
rect 4672 10656 4678 10668
rect 5184 10665 5212 10764
rect 5442 10752 5448 10764
rect 5500 10752 5506 10804
rect 5629 10795 5687 10801
rect 5629 10761 5641 10795
rect 5675 10792 5687 10795
rect 7834 10792 7840 10804
rect 5675 10764 7696 10792
rect 7795 10764 7840 10792
rect 5675 10761 5687 10764
rect 5629 10755 5687 10761
rect 6086 10684 6092 10736
rect 6144 10724 6150 10736
rect 7668 10724 7696 10764
rect 7834 10752 7840 10764
rect 7892 10752 7898 10804
rect 6144 10696 6500 10724
rect 7668 10696 7788 10724
rect 6144 10684 6150 10696
rect 4893 10659 4951 10665
rect 4893 10656 4905 10659
rect 4672 10628 4905 10656
rect 4672 10616 4678 10628
rect 4893 10625 4905 10628
rect 4939 10625 4951 10659
rect 4893 10619 4951 10625
rect 5169 10659 5227 10665
rect 5169 10625 5181 10659
rect 5215 10625 5227 10659
rect 5169 10619 5227 10625
rect 5534 10616 5540 10668
rect 5592 10656 5598 10668
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5592 10628 6009 10656
rect 5592 10616 5598 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 6178 10656 6184 10668
rect 6139 10628 6184 10656
rect 5997 10619 6055 10625
rect 6178 10616 6184 10628
rect 6236 10616 6242 10668
rect 6472 10656 6500 10696
rect 6472 10628 6684 10656
rect 1305 10591 1363 10597
rect 1305 10557 1317 10591
rect 1351 10588 1363 10591
rect 1854 10588 1860 10600
rect 1351 10560 1860 10588
rect 1351 10557 1363 10560
rect 1305 10551 1363 10557
rect 1854 10548 1860 10560
rect 1912 10548 1918 10600
rect 2130 10588 2136 10600
rect 2091 10560 2136 10588
rect 2130 10548 2136 10560
rect 2188 10548 2194 10600
rect 4169 10591 4227 10597
rect 4169 10557 4181 10591
rect 4215 10588 4227 10591
rect 6656 10588 6684 10628
rect 6730 10616 6736 10668
rect 6788 10656 6794 10668
rect 6917 10659 6975 10665
rect 6917 10656 6929 10659
rect 6788 10628 6929 10656
rect 6788 10616 6794 10628
rect 6917 10625 6929 10628
rect 6963 10625 6975 10659
rect 6917 10619 6975 10625
rect 7101 10659 7159 10665
rect 7101 10625 7113 10659
rect 7147 10656 7159 10659
rect 7190 10656 7196 10668
rect 7147 10628 7196 10656
rect 7147 10625 7159 10628
rect 7101 10619 7159 10625
rect 7190 10616 7196 10628
rect 7248 10616 7254 10668
rect 7653 10659 7711 10665
rect 7653 10625 7665 10659
rect 7699 10658 7711 10659
rect 7760 10658 7788 10696
rect 7699 10630 7788 10658
rect 7929 10659 7987 10665
rect 7699 10625 7711 10630
rect 7653 10619 7711 10625
rect 7929 10625 7941 10659
rect 7975 10656 7987 10659
rect 8110 10656 8116 10668
rect 7975 10628 8116 10656
rect 7975 10625 7987 10628
rect 7929 10619 7987 10625
rect 8110 10616 8116 10628
rect 8168 10616 8174 10668
rect 8297 10659 8355 10665
rect 8297 10625 8309 10659
rect 8343 10625 8355 10659
rect 9306 10656 9312 10668
rect 9267 10628 9312 10656
rect 8297 10619 8355 10625
rect 8312 10588 8340 10619
rect 9306 10616 9312 10628
rect 9364 10616 9370 10668
rect 4215 10560 6408 10588
rect 6656 10560 8340 10588
rect 4215 10557 4227 10560
rect 4169 10551 4227 10557
rect 5276 10492 5948 10520
rect 4798 10452 4804 10464
rect 4759 10424 4804 10452
rect 4798 10412 4804 10424
rect 4856 10452 4862 10464
rect 5276 10461 5304 10492
rect 5261 10455 5319 10461
rect 5261 10452 5273 10455
rect 4856 10424 5273 10452
rect 4856 10412 4862 10424
rect 5261 10421 5273 10424
rect 5307 10421 5319 10455
rect 5810 10452 5816 10464
rect 5771 10424 5816 10452
rect 5261 10415 5319 10421
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 5920 10452 5948 10492
rect 6273 10455 6331 10461
rect 6273 10452 6285 10455
rect 5920 10424 6285 10452
rect 6273 10421 6285 10424
rect 6319 10421 6331 10455
rect 6380 10452 6408 10560
rect 8386 10548 8392 10600
rect 8444 10588 8450 10600
rect 9401 10591 9459 10597
rect 9401 10588 9413 10591
rect 8444 10560 9413 10588
rect 8444 10548 8450 10560
rect 9401 10557 9413 10560
rect 9447 10557 9459 10591
rect 9401 10551 9459 10557
rect 6641 10523 6699 10529
rect 6641 10489 6653 10523
rect 6687 10520 6699 10523
rect 7558 10520 7564 10532
rect 6687 10492 7564 10520
rect 6687 10489 6699 10492
rect 6641 10483 6699 10489
rect 7558 10480 7564 10492
rect 7616 10480 7622 10532
rect 8481 10523 8539 10529
rect 8481 10489 8493 10523
rect 8527 10520 8539 10523
rect 8527 10492 16574 10520
rect 8527 10489 8539 10492
rect 8481 10483 8539 10489
rect 16546 10464 16574 10492
rect 7098 10452 7104 10464
rect 6380 10424 7104 10452
rect 6273 10415 6331 10421
rect 7098 10412 7104 10424
rect 7156 10412 7162 10464
rect 7282 10452 7288 10464
rect 7243 10424 7288 10452
rect 7282 10412 7288 10424
rect 7340 10412 7346 10464
rect 7466 10452 7472 10464
rect 7427 10424 7472 10452
rect 7466 10412 7472 10424
rect 7524 10412 7530 10464
rect 8110 10452 8116 10464
rect 8071 10424 8116 10452
rect 8110 10412 8116 10424
rect 8168 10412 8174 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 8665 10455 8723 10461
rect 8665 10452 8677 10455
rect 8352 10424 8677 10452
rect 8352 10412 8358 10424
rect 8665 10421 8677 10424
rect 8711 10421 8723 10455
rect 16546 10424 16580 10464
rect 8665 10415 8723 10421
rect 16574 10412 16580 10424
rect 16632 10412 16638 10464
rect 920 10362 9844 10384
rect 920 10310 2566 10362
rect 2618 10310 2630 10362
rect 2682 10310 2694 10362
rect 2746 10310 2758 10362
rect 2810 10310 2822 10362
rect 2874 10310 7566 10362
rect 7618 10310 7630 10362
rect 7682 10310 7694 10362
rect 7746 10310 7758 10362
rect 7810 10310 7822 10362
rect 7874 10310 9844 10362
rect 920 10288 9844 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 4433 10251 4491 10257
rect 4433 10248 4445 10251
rect 1544 10220 4445 10248
rect 1544 10208 1550 10220
rect 4433 10217 4445 10220
rect 4479 10248 4491 10251
rect 6730 10248 6736 10260
rect 4479 10220 6736 10248
rect 4479 10217 4491 10220
rect 4433 10211 4491 10217
rect 6730 10208 6736 10220
rect 6788 10208 6794 10260
rect 7190 10208 7196 10260
rect 7248 10248 7254 10260
rect 8757 10251 8815 10257
rect 8757 10248 8769 10251
rect 7248 10220 8769 10248
rect 7248 10208 7254 10220
rect 8757 10217 8769 10220
rect 8803 10217 8815 10251
rect 8757 10211 8815 10217
rect 2130 10140 2136 10192
rect 2188 10180 2194 10192
rect 2685 10183 2743 10189
rect 2685 10180 2697 10183
rect 2188 10152 2697 10180
rect 2188 10140 2194 10152
rect 2685 10149 2697 10152
rect 2731 10149 2743 10183
rect 2685 10143 2743 10149
rect 3234 10140 3240 10192
rect 3292 10180 3298 10192
rect 3605 10183 3663 10189
rect 3605 10180 3617 10183
rect 3292 10152 3617 10180
rect 3292 10140 3298 10152
rect 3605 10149 3617 10152
rect 3651 10149 3663 10183
rect 3605 10143 3663 10149
rect 8202 10140 8208 10192
rect 8260 10180 8266 10192
rect 8481 10183 8539 10189
rect 8481 10180 8493 10183
rect 8260 10152 8493 10180
rect 8260 10140 8266 10152
rect 8481 10149 8493 10152
rect 8527 10149 8539 10183
rect 8481 10143 8539 10149
rect 1305 10115 1363 10121
rect 1305 10081 1317 10115
rect 1351 10112 1363 10115
rect 1351 10084 2084 10112
rect 1351 10081 1363 10084
rect 1305 10075 1363 10081
rect 2056 10053 2084 10084
rect 7282 10072 7288 10124
rect 7340 10112 7346 10124
rect 8297 10115 8355 10121
rect 8297 10112 8309 10115
rect 7340 10084 8309 10112
rect 7340 10072 7346 10084
rect 8297 10081 8309 10084
rect 8343 10081 8355 10115
rect 9490 10112 9496 10124
rect 8297 10075 8355 10081
rect 8588 10084 9496 10112
rect 1949 10047 2007 10053
rect 1949 10013 1961 10047
rect 1995 10013 2007 10047
rect 1949 10007 2007 10013
rect 2041 10047 2099 10053
rect 2041 10013 2053 10047
rect 2087 10013 2099 10047
rect 2041 10007 2099 10013
rect 1964 9976 1992 10007
rect 3050 10004 3056 10056
rect 3108 10044 3114 10056
rect 3421 10047 3479 10053
rect 3421 10044 3433 10047
rect 3108 10016 3433 10044
rect 3108 10004 3114 10016
rect 3421 10013 3433 10016
rect 3467 10013 3479 10047
rect 3786 10044 3792 10056
rect 3747 10016 3792 10044
rect 3421 10007 3479 10013
rect 3786 10004 3792 10016
rect 3844 10004 3850 10056
rect 4890 10004 4896 10056
rect 4948 10044 4954 10056
rect 5721 10047 5779 10053
rect 5721 10044 5733 10047
rect 4948 10016 5733 10044
rect 4948 10004 4954 10016
rect 5721 10013 5733 10016
rect 5767 10013 5779 10047
rect 5721 10007 5779 10013
rect 6178 10004 6184 10056
rect 6236 10044 6242 10056
rect 6457 10047 6515 10053
rect 6457 10044 6469 10047
rect 6236 10016 6469 10044
rect 6236 10004 6242 10016
rect 6457 10013 6469 10016
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 7929 10047 7987 10053
rect 7929 10013 7941 10047
rect 7975 10044 7987 10047
rect 8478 10044 8484 10056
rect 7975 10016 8484 10044
rect 7975 10013 7987 10016
rect 7929 10007 7987 10013
rect 8478 10004 8484 10016
rect 8536 10004 8542 10056
rect 8588 10053 8616 10084
rect 9490 10072 9496 10084
rect 9548 10072 9554 10124
rect 8573 10047 8631 10053
rect 8573 10013 8585 10047
rect 8619 10013 8631 10047
rect 9398 10044 9404 10056
rect 9359 10016 9404 10044
rect 8573 10007 8631 10013
rect 9398 10004 9404 10016
rect 9456 10004 9462 10056
rect 2777 9979 2835 9985
rect 2777 9976 2789 9979
rect 1964 9948 2789 9976
rect 2777 9945 2789 9948
rect 2823 9945 2835 9979
rect 2777 9939 2835 9945
rect 7466 9936 7472 9988
rect 7524 9936 7530 9988
rect 8412 9948 16574 9976
rect 5897 9911 5955 9917
rect 5897 9877 5909 9911
rect 5943 9908 5955 9911
rect 8412 9908 8440 9948
rect 5943 9880 8440 9908
rect 5943 9877 5955 9880
rect 5897 9871 5955 9877
rect 920 9818 9844 9840
rect 920 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 5194 9818
rect 5246 9766 5258 9818
rect 5310 9766 5322 9818
rect 5374 9766 9844 9818
rect 920 9744 9844 9766
rect 1854 9664 1860 9716
rect 1912 9664 1918 9716
rect 7282 9664 7288 9716
rect 7340 9704 7346 9716
rect 8202 9704 8208 9716
rect 7340 9676 8208 9704
rect 7340 9664 7346 9676
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 9490 9704 9496 9716
rect 9451 9676 9496 9704
rect 9490 9664 9496 9676
rect 9548 9664 9554 9716
rect 16546 9704 16574 9948
rect 16666 9704 16672 9716
rect 16546 9676 16672 9704
rect 16666 9664 16672 9676
rect 16724 9664 16730 9716
rect 1486 9636 1492 9648
rect 1447 9608 1492 9636
rect 1486 9596 1492 9608
rect 1544 9596 1550 9648
rect 1872 9636 1900 9664
rect 1872 9608 1978 9636
rect 4522 9596 4528 9648
rect 4580 9596 4586 9648
rect 7926 9596 7932 9648
rect 7984 9596 7990 9648
rect 3142 9528 3148 9580
rect 3200 9568 3206 9580
rect 3329 9571 3387 9577
rect 3329 9568 3341 9571
rect 3200 9540 3341 9568
rect 3200 9528 3206 9540
rect 3329 9537 3341 9540
rect 3375 9537 3387 9571
rect 3329 9531 3387 9537
rect 3418 9528 3424 9580
rect 3476 9568 3482 9580
rect 5261 9571 5319 9577
rect 3476 9540 3521 9568
rect 3476 9528 3482 9540
rect 5261 9537 5273 9571
rect 5307 9568 5319 9571
rect 5810 9568 5816 9580
rect 5307 9540 5816 9568
rect 5307 9537 5319 9540
rect 5261 9531 5319 9537
rect 5810 9528 5816 9540
rect 5868 9528 5874 9580
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 6365 9571 6423 9577
rect 6365 9568 6377 9571
rect 6328 9540 6377 9568
rect 6328 9528 6334 9540
rect 6365 9537 6377 9540
rect 6411 9537 6423 9571
rect 6546 9568 6552 9580
rect 6507 9540 6552 9568
rect 6365 9531 6423 9537
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 6825 9571 6883 9577
rect 6825 9537 6837 9571
rect 6871 9568 6883 9571
rect 7006 9568 7012 9580
rect 6871 9540 7012 9568
rect 6871 9537 6883 9540
rect 6825 9531 6883 9537
rect 7006 9528 7012 9540
rect 7064 9528 7070 9580
rect 8110 9528 8116 9580
rect 8168 9568 8174 9580
rect 8665 9571 8723 9577
rect 8665 9568 8677 9571
rect 8168 9540 8677 9568
rect 8168 9528 8174 9540
rect 8665 9537 8677 9540
rect 8711 9537 8723 9571
rect 8665 9531 8723 9537
rect 1213 9503 1271 9509
rect 1213 9469 1225 9503
rect 1259 9500 1271 9503
rect 3789 9503 3847 9509
rect 1259 9472 2774 9500
rect 1259 9469 1271 9472
rect 1213 9463 1271 9469
rect 2746 9432 2774 9472
rect 3789 9469 3801 9503
rect 3835 9500 3847 9503
rect 4062 9500 4068 9512
rect 3835 9472 4068 9500
rect 3835 9469 3847 9472
rect 3789 9463 3847 9469
rect 4062 9460 4068 9472
rect 4120 9460 4126 9512
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 6454 9500 6460 9512
rect 5408 9472 6460 9500
rect 5408 9460 5414 9472
rect 6454 9460 6460 9472
rect 6512 9460 6518 9512
rect 7193 9503 7251 9509
rect 7193 9500 7205 9503
rect 6932 9472 7205 9500
rect 3418 9432 3424 9444
rect 2746 9404 3424 9432
rect 3418 9392 3424 9404
rect 3476 9392 3482 9444
rect 6086 9432 6092 9444
rect 5184 9404 6092 9432
rect 2961 9367 3019 9373
rect 2961 9333 2973 9367
rect 3007 9364 3019 9367
rect 3050 9364 3056 9376
rect 3007 9336 3056 9364
rect 3007 9333 3019 9336
rect 2961 9327 3019 9333
rect 3050 9324 3056 9336
rect 3108 9324 3114 9376
rect 3145 9367 3203 9373
rect 3145 9333 3157 9367
rect 3191 9364 3203 9367
rect 3234 9364 3240 9376
rect 3191 9336 3240 9364
rect 3191 9333 3203 9336
rect 3145 9327 3203 9333
rect 3234 9324 3240 9336
rect 3292 9324 3298 9376
rect 4154 9324 4160 9376
rect 4212 9364 4218 9376
rect 5184 9364 5212 9404
rect 6086 9392 6092 9404
rect 6144 9432 6150 9444
rect 6181 9435 6239 9441
rect 6181 9432 6193 9435
rect 6144 9404 6193 9432
rect 6144 9392 6150 9404
rect 6181 9401 6193 9404
rect 6227 9401 6239 9435
rect 6730 9432 6736 9444
rect 6691 9404 6736 9432
rect 6181 9395 6239 9401
rect 6730 9392 6736 9404
rect 6788 9392 6794 9444
rect 4212 9336 5212 9364
rect 5825 9367 5883 9373
rect 4212 9324 4218 9336
rect 5825 9333 5837 9367
rect 5871 9364 5883 9367
rect 6822 9364 6828 9376
rect 5871 9336 6828 9364
rect 5871 9333 5883 9336
rect 5825 9327 5883 9333
rect 6822 9324 6828 9336
rect 6880 9324 6886 9376
rect 6932 9364 6960 9472
rect 7193 9469 7205 9472
rect 7239 9469 7251 9503
rect 7193 9463 7251 9469
rect 8294 9364 8300 9376
rect 6932 9336 8300 9364
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 9214 9364 9220 9376
rect 9272 9373 9278 9376
rect 9183 9336 9220 9364
rect 9214 9324 9220 9336
rect 9272 9327 9283 9373
rect 9272 9324 9278 9327
rect 920 9274 9844 9296
rect 920 9222 2566 9274
rect 2618 9222 2630 9274
rect 2682 9222 2694 9274
rect 2746 9222 2758 9274
rect 2810 9222 2822 9274
rect 2874 9222 7566 9274
rect 7618 9222 7630 9274
rect 7682 9222 7694 9274
rect 7746 9222 7758 9274
rect 7810 9222 7822 9274
rect 7874 9222 9844 9274
rect 920 9200 9844 9222
rect 1394 9120 1400 9172
rect 1452 9160 1458 9172
rect 1673 9163 1731 9169
rect 1673 9160 1685 9163
rect 1452 9132 1685 9160
rect 1452 9120 1458 9132
rect 1504 9024 1532 9132
rect 1673 9129 1685 9132
rect 1719 9129 1731 9163
rect 1673 9123 1731 9129
rect 2317 9163 2375 9169
rect 2317 9129 2329 9163
rect 2363 9160 2375 9163
rect 2406 9160 2412 9172
rect 2363 9132 2412 9160
rect 2363 9129 2375 9132
rect 2317 9123 2375 9129
rect 2406 9120 2412 9132
rect 2464 9160 2470 9172
rect 2777 9163 2835 9169
rect 2777 9160 2789 9163
rect 2464 9132 2789 9160
rect 2464 9120 2470 9132
rect 2777 9129 2789 9132
rect 2823 9129 2835 9163
rect 3142 9160 3148 9172
rect 3103 9132 3148 9160
rect 2777 9123 2835 9129
rect 3142 9120 3148 9132
rect 3200 9120 3206 9172
rect 3973 9163 4031 9169
rect 3973 9129 3985 9163
rect 4019 9160 4031 9163
rect 5350 9160 5356 9172
rect 4019 9132 5356 9160
rect 4019 9129 4031 9132
rect 3973 9123 4031 9129
rect 1578 9052 1584 9104
rect 1636 9092 1642 9104
rect 3988 9092 4016 9123
rect 5350 9120 5356 9132
rect 5408 9160 5414 9172
rect 5994 9160 6000 9172
rect 5408 9132 6000 9160
rect 5408 9120 5414 9132
rect 5994 9120 6000 9132
rect 6052 9120 6058 9172
rect 6546 9120 6552 9172
rect 6604 9160 6610 9172
rect 8846 9160 8852 9172
rect 6604 9132 8852 9160
rect 6604 9120 6610 9132
rect 8846 9120 8852 9132
rect 8904 9120 8910 9172
rect 9398 9160 9404 9172
rect 9359 9132 9404 9160
rect 9398 9120 9404 9132
rect 9456 9120 9462 9172
rect 1636 9064 4016 9092
rect 4893 9095 4951 9101
rect 1636 9052 1642 9064
rect 4893 9061 4905 9095
rect 4939 9092 4951 9095
rect 5166 9092 5172 9104
rect 4939 9064 5172 9092
rect 4939 9061 4951 9064
rect 4893 9055 4951 9061
rect 5166 9052 5172 9064
rect 5224 9052 5230 9104
rect 5261 9095 5319 9101
rect 5261 9061 5273 9095
rect 5307 9061 5319 9095
rect 5718 9092 5724 9104
rect 5679 9064 5724 9092
rect 5261 9055 5319 9061
rect 2501 9027 2559 9033
rect 1504 8996 2084 9024
rect 1486 8956 1492 8968
rect 1447 8928 1492 8956
rect 1486 8916 1492 8928
rect 1544 8916 1550 8968
rect 1670 8916 1676 8968
rect 1728 8956 1734 8968
rect 2056 8965 2084 8996
rect 2501 8993 2513 9027
rect 2547 9024 2559 9027
rect 3786 9024 3792 9036
rect 2547 8996 3792 9024
rect 2547 8993 2559 8996
rect 2501 8987 2559 8993
rect 3786 8984 3792 8996
rect 3844 8984 3850 9036
rect 4798 9024 4804 9036
rect 3988 8996 4804 9024
rect 1949 8959 2007 8965
rect 1949 8956 1961 8959
rect 1728 8928 1961 8956
rect 1728 8916 1734 8928
rect 1949 8925 1961 8928
rect 1995 8925 2007 8959
rect 1949 8919 2007 8925
rect 2041 8959 2099 8965
rect 2041 8925 2053 8959
rect 2087 8925 2099 8959
rect 2041 8919 2099 8925
rect 2685 8959 2743 8965
rect 2685 8925 2697 8959
rect 2731 8956 2743 8959
rect 2731 8928 3004 8956
rect 2731 8925 2743 8928
rect 2685 8919 2743 8925
rect 1305 8891 1363 8897
rect 1305 8857 1317 8891
rect 1351 8888 1363 8891
rect 1394 8888 1400 8900
rect 1351 8860 1400 8888
rect 1351 8857 1363 8860
rect 1305 8851 1363 8857
rect 1394 8848 1400 8860
rect 1452 8888 1458 8900
rect 1452 8860 1992 8888
rect 1452 8848 1458 8860
rect 1964 8832 1992 8860
rect 2406 8848 2412 8900
rect 2464 8888 2470 8900
rect 2976 8888 3004 8928
rect 3326 8916 3332 8968
rect 3384 8956 3390 8968
rect 3605 8959 3663 8965
rect 3605 8956 3617 8959
rect 3384 8928 3617 8956
rect 3384 8916 3390 8928
rect 3605 8925 3617 8928
rect 3651 8925 3663 8959
rect 3605 8919 3663 8925
rect 3421 8891 3479 8897
rect 3421 8888 3433 8891
rect 2464 8860 2774 8888
rect 2976 8860 3433 8888
rect 2464 8848 2470 8860
rect 1762 8780 1768 8832
rect 1820 8820 1826 8832
rect 1857 8823 1915 8829
rect 1857 8820 1869 8823
rect 1820 8792 1869 8820
rect 1820 8780 1826 8792
rect 1857 8789 1869 8792
rect 1903 8789 1915 8823
rect 1857 8783 1915 8789
rect 1946 8780 1952 8832
rect 2004 8780 2010 8832
rect 2746 8820 2774 8860
rect 3421 8857 3433 8860
rect 3467 8888 3479 8891
rect 3510 8888 3516 8900
rect 3467 8860 3516 8888
rect 3467 8857 3479 8860
rect 3421 8851 3479 8857
rect 3510 8848 3516 8860
rect 3568 8848 3574 8900
rect 3988 8888 4016 8996
rect 4798 8984 4804 8996
rect 4856 9024 4862 9036
rect 5276 9024 5304 9055
rect 5718 9052 5724 9064
rect 5776 9052 5782 9104
rect 6089 9095 6147 9101
rect 6089 9061 6101 9095
rect 6135 9092 6147 9095
rect 6178 9092 6184 9104
rect 6135 9064 6184 9092
rect 6135 9061 6147 9064
rect 6089 9055 6147 9061
rect 6178 9052 6184 9064
rect 6236 9052 6242 9104
rect 4856 8996 5304 9024
rect 5368 8996 6224 9024
rect 4856 8984 4862 8996
rect 4246 8956 4252 8968
rect 4207 8928 4252 8956
rect 4246 8916 4252 8928
rect 4304 8916 4310 8968
rect 4525 8959 4583 8965
rect 4525 8925 4537 8959
rect 4571 8956 4583 8959
rect 4614 8956 4620 8968
rect 4571 8928 4620 8956
rect 4571 8925 4583 8928
rect 4525 8919 4583 8925
rect 4614 8916 4620 8928
rect 4672 8916 4678 8968
rect 4982 8916 4988 8968
rect 5040 8956 5046 8968
rect 5169 8959 5227 8965
rect 5169 8956 5181 8959
rect 5040 8928 5181 8956
rect 5040 8916 5046 8928
rect 5169 8925 5181 8928
rect 5215 8956 5227 8959
rect 5368 8956 5396 8996
rect 5215 8928 5396 8956
rect 5445 8959 5503 8965
rect 5215 8925 5227 8928
rect 5169 8919 5227 8925
rect 5445 8925 5457 8959
rect 5491 8956 5503 8959
rect 5534 8956 5540 8968
rect 5491 8928 5540 8956
rect 5491 8925 5503 8928
rect 5445 8919 5503 8925
rect 5534 8916 5540 8928
rect 5592 8916 5598 8968
rect 5902 8956 5908 8968
rect 5863 8928 5908 8956
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 6196 8900 6224 8996
rect 6362 8984 6368 9036
rect 6420 9024 6426 9036
rect 8021 9027 8079 9033
rect 8021 9024 8033 9027
rect 6420 8996 8033 9024
rect 6420 8984 6426 8996
rect 8021 8993 8033 8996
rect 8067 8993 8079 9027
rect 8021 8987 8079 8993
rect 8036 8956 8064 8987
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 9122 9024 9128 9036
rect 8444 8996 9128 9024
rect 8444 8984 8450 8996
rect 9122 8984 9128 8996
rect 9180 8984 9186 9036
rect 8297 8959 8355 8965
rect 8297 8956 8309 8959
rect 8036 8928 8309 8956
rect 8297 8925 8309 8928
rect 8343 8956 8355 8959
rect 8570 8956 8576 8968
rect 8343 8928 8576 8956
rect 8343 8925 8355 8928
rect 8297 8919 8355 8925
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 8754 8956 8760 8968
rect 8715 8928 8760 8956
rect 8754 8916 8760 8928
rect 8812 8916 8818 8968
rect 3620 8860 4016 8888
rect 4065 8891 4123 8897
rect 3620 8820 3648 8860
rect 4065 8857 4077 8891
rect 4111 8888 4123 8891
rect 4338 8888 4344 8900
rect 4111 8860 4344 8888
rect 4111 8857 4123 8860
rect 4065 8851 4123 8857
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 4709 8891 4767 8897
rect 4709 8857 4721 8891
rect 4755 8888 4767 8891
rect 5718 8888 5724 8900
rect 4755 8860 5724 8888
rect 4755 8857 4767 8860
rect 4709 8851 4767 8857
rect 5718 8848 5724 8860
rect 5776 8848 5782 8900
rect 6178 8888 6184 8900
rect 6091 8860 6184 8888
rect 6178 8848 6184 8860
rect 6236 8888 6242 8900
rect 7745 8891 7803 8897
rect 6236 8860 6578 8888
rect 6236 8848 6242 8860
rect 7745 8857 7757 8891
rect 7791 8888 7803 8891
rect 7834 8888 7840 8900
rect 7791 8860 7840 8888
rect 7791 8857 7803 8860
rect 7745 8851 7803 8857
rect 7834 8848 7840 8860
rect 7892 8848 7898 8900
rect 8386 8888 8392 8900
rect 8036 8860 8392 8888
rect 3786 8820 3792 8832
rect 2746 8792 3648 8820
rect 3747 8792 3792 8820
rect 3786 8780 3792 8792
rect 3844 8780 3850 8832
rect 4433 8823 4491 8829
rect 4433 8789 4445 8823
rect 4479 8820 4491 8823
rect 4798 8820 4804 8832
rect 4479 8792 4804 8820
rect 4479 8789 4491 8792
rect 4433 8783 4491 8789
rect 4798 8780 4804 8792
rect 4856 8780 4862 8832
rect 4985 8823 5043 8829
rect 4985 8789 4997 8823
rect 5031 8820 5043 8823
rect 5442 8820 5448 8832
rect 5031 8792 5448 8820
rect 5031 8789 5043 8792
rect 4985 8783 5043 8789
rect 5442 8780 5448 8792
rect 5500 8780 5506 8832
rect 6273 8823 6331 8829
rect 6273 8789 6285 8823
rect 6319 8820 6331 8823
rect 8036 8820 8064 8860
rect 8386 8848 8392 8860
rect 8444 8848 8450 8900
rect 8496 8860 16574 8888
rect 6319 8792 8064 8820
rect 8205 8823 8263 8829
rect 6319 8789 6331 8792
rect 6273 8783 6331 8789
rect 8205 8789 8217 8823
rect 8251 8820 8263 8823
rect 8294 8820 8300 8832
rect 8251 8792 8300 8820
rect 8251 8789 8263 8792
rect 8205 8783 8263 8789
rect 8294 8780 8300 8792
rect 8352 8780 8358 8832
rect 8496 8829 8524 8860
rect 16546 8832 16574 8860
rect 8481 8823 8539 8829
rect 8481 8789 8493 8823
rect 8527 8789 8539 8823
rect 16546 8792 16580 8832
rect 8481 8783 8539 8789
rect 16574 8780 16580 8792
rect 16632 8780 16638 8832
rect 920 8730 9844 8752
rect 920 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 5194 8730
rect 5246 8678 5258 8730
rect 5310 8678 5322 8730
rect 5374 8678 9844 8730
rect 920 8656 9844 8678
rect 1581 8619 1639 8625
rect 1581 8585 1593 8619
rect 1627 8616 1639 8619
rect 3142 8616 3148 8628
rect 1627 8588 3148 8616
rect 1627 8585 1639 8588
rect 1581 8579 1639 8585
rect 3142 8576 3148 8588
rect 3200 8576 3206 8628
rect 5534 8616 5540 8628
rect 4172 8588 5540 8616
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 1578 8440 1584 8492
rect 1636 8480 1642 8492
rect 1673 8483 1731 8489
rect 1673 8480 1685 8483
rect 1636 8452 1685 8480
rect 1636 8440 1642 8452
rect 1673 8449 1685 8452
rect 1719 8449 1731 8483
rect 1673 8443 1731 8449
rect 1762 8440 1768 8492
rect 1820 8480 1826 8492
rect 3605 8483 3663 8489
rect 1820 8452 1865 8480
rect 1820 8440 1826 8452
rect 3605 8449 3617 8483
rect 3651 8480 3663 8483
rect 3786 8480 3792 8492
rect 3651 8452 3792 8480
rect 3651 8449 3663 8452
rect 3605 8443 3663 8449
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 4172 8480 4200 8588
rect 5534 8576 5540 8588
rect 5592 8616 5598 8628
rect 5997 8619 6055 8625
rect 5592 8588 5856 8616
rect 5592 8576 5598 8588
rect 4246 8508 4252 8560
rect 4304 8548 4310 8560
rect 5445 8551 5503 8557
rect 5445 8548 5457 8551
rect 4304 8520 5457 8548
rect 4304 8508 4310 8520
rect 5445 8517 5457 8520
rect 5491 8517 5503 8551
rect 5445 8511 5503 8517
rect 5629 8551 5687 8557
rect 5629 8517 5641 8551
rect 5675 8548 5687 8551
rect 5718 8548 5724 8560
rect 5675 8520 5724 8548
rect 5675 8517 5687 8520
rect 5629 8511 5687 8517
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 4172 8452 4353 8480
rect 1397 8415 1455 8421
rect 1397 8381 1409 8415
rect 1443 8412 1455 8415
rect 1854 8412 1860 8424
rect 1443 8384 1860 8412
rect 1443 8381 1455 8384
rect 1397 8375 1455 8381
rect 1854 8372 1860 8384
rect 1912 8372 1918 8424
rect 2130 8412 2136 8424
rect 2091 8384 2136 8412
rect 2130 8372 2136 8384
rect 2188 8372 2194 8424
rect 1872 8276 1900 8372
rect 4172 8344 4200 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4341 8443 4399 8449
rect 4430 8440 4436 8492
rect 4488 8480 4494 8492
rect 4982 8480 4988 8492
rect 4488 8452 4988 8480
rect 4488 8440 4494 8452
rect 4982 8440 4988 8452
rect 5040 8440 5046 8492
rect 5169 8483 5227 8489
rect 5169 8449 5181 8483
rect 5215 8480 5227 8483
rect 5644 8480 5672 8511
rect 5718 8508 5724 8520
rect 5776 8508 5782 8560
rect 5828 8557 5856 8588
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6178 8616 6184 8628
rect 6043 8588 6184 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6178 8576 6184 8588
rect 6236 8576 6242 8628
rect 7193 8619 7251 8625
rect 7193 8585 7205 8619
rect 7239 8616 7251 8619
rect 8754 8616 8760 8628
rect 7239 8588 8760 8616
rect 7239 8585 7251 8588
rect 7193 8579 7251 8585
rect 8754 8576 8760 8588
rect 8812 8576 8818 8628
rect 9122 8576 9128 8628
rect 9180 8616 9186 8628
rect 9401 8619 9459 8625
rect 9180 8588 9260 8616
rect 9180 8576 9186 8588
rect 5813 8551 5871 8557
rect 5813 8517 5825 8551
rect 5859 8517 5871 8551
rect 6196 8548 6224 8576
rect 7466 8548 7472 8560
rect 6196 8520 7472 8548
rect 5813 8511 5871 8517
rect 7466 8508 7472 8520
rect 7524 8548 7530 8560
rect 7524 8534 7682 8548
rect 7524 8520 7696 8534
rect 7524 8508 7530 8520
rect 5215 8452 5672 8480
rect 5215 8449 5227 8452
rect 5169 8443 5227 8449
rect 5902 8440 5908 8492
rect 5960 8480 5966 8492
rect 6273 8483 6331 8489
rect 6273 8480 6285 8483
rect 5960 8452 6285 8480
rect 5960 8440 5966 8452
rect 6273 8449 6285 8452
rect 6319 8449 6331 8483
rect 6273 8443 6331 8449
rect 6549 8483 6607 8489
rect 6549 8449 6561 8483
rect 6595 8449 6607 8483
rect 6549 8443 6607 8449
rect 4801 8415 4859 8421
rect 4801 8381 4813 8415
rect 4847 8412 4859 8415
rect 6178 8412 6184 8424
rect 4847 8384 6184 8412
rect 4847 8381 4859 8384
rect 4801 8375 4859 8381
rect 6178 8372 6184 8384
rect 6236 8372 6242 8424
rect 6454 8372 6460 8424
rect 6512 8412 6518 8424
rect 6564 8412 6592 8443
rect 7377 8415 7435 8421
rect 7377 8412 7389 8415
rect 6512 8384 7389 8412
rect 6512 8372 6518 8384
rect 7377 8381 7389 8384
rect 7423 8381 7435 8415
rect 7668 8412 7696 8520
rect 8570 8508 8576 8560
rect 8628 8548 8634 8560
rect 8628 8520 9168 8548
rect 8628 8508 8634 8520
rect 9140 8489 9168 8520
rect 9232 8489 9260 8588
rect 9401 8585 9413 8619
rect 9447 8616 9459 8619
rect 16574 8616 16580 8628
rect 9447 8588 16580 8616
rect 9447 8585 9459 8588
rect 9401 8579 9459 8585
rect 16574 8576 16580 8588
rect 16632 8576 16638 8628
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 9125 8443 9183 8449
rect 9217 8483 9275 8489
rect 9217 8449 9229 8483
rect 9263 8449 9275 8483
rect 9217 8443 9275 8449
rect 8202 8412 8208 8424
rect 7668 8384 8208 8412
rect 7377 8375 7435 8381
rect 8202 8372 8208 8384
rect 8260 8372 8266 8424
rect 8386 8372 8392 8424
rect 8444 8412 8450 8424
rect 8754 8412 8760 8424
rect 8444 8384 8760 8412
rect 8444 8372 8450 8384
rect 8754 8372 8760 8384
rect 8812 8412 8818 8424
rect 8849 8415 8907 8421
rect 8849 8412 8861 8415
rect 8812 8384 8861 8412
rect 8812 8372 8818 8384
rect 8849 8381 8861 8384
rect 8895 8381 8907 8415
rect 8849 8375 8907 8381
rect 5353 8347 5411 8353
rect 3068 8316 4200 8344
rect 4448 8316 5304 8344
rect 3068 8276 3096 8316
rect 1872 8248 3096 8276
rect 4169 8279 4227 8285
rect 4169 8245 4181 8279
rect 4215 8276 4227 8279
rect 4448 8276 4476 8316
rect 4614 8276 4620 8288
rect 4215 8248 4476 8276
rect 4575 8248 4620 8276
rect 4215 8245 4227 8248
rect 4169 8239 4227 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 5276 8276 5304 8316
rect 5353 8313 5365 8347
rect 5399 8344 5411 8347
rect 5810 8344 5816 8356
rect 5399 8316 5816 8344
rect 5399 8313 5411 8316
rect 5353 8307 5411 8313
rect 5810 8304 5816 8316
rect 5868 8304 5874 8356
rect 6822 8304 6828 8356
rect 6880 8344 6886 8356
rect 6880 8316 7880 8344
rect 6880 8304 6886 8316
rect 5442 8276 5448 8288
rect 5276 8248 5448 8276
rect 5442 8236 5448 8248
rect 5500 8236 5506 8288
rect 6362 8276 6368 8288
rect 6323 8248 6368 8276
rect 6362 8236 6368 8248
rect 6420 8236 6426 8288
rect 7006 8236 7012 8288
rect 7064 8276 7070 8288
rect 7190 8276 7196 8288
rect 7064 8248 7196 8276
rect 7064 8236 7070 8248
rect 7190 8236 7196 8248
rect 7248 8236 7254 8288
rect 7852 8276 7880 8316
rect 9030 8276 9036 8288
rect 7852 8248 9036 8276
rect 9030 8236 9036 8248
rect 9088 8236 9094 8288
rect 920 8186 9844 8208
rect 920 8134 2566 8186
rect 2618 8134 2630 8186
rect 2682 8134 2694 8186
rect 2746 8134 2758 8186
rect 2810 8134 2822 8186
rect 2874 8134 7566 8186
rect 7618 8134 7630 8186
rect 7682 8134 7694 8186
rect 7746 8134 7758 8186
rect 7810 8134 7822 8186
rect 7874 8134 9844 8186
rect 920 8112 9844 8134
rect 2130 8032 2136 8084
rect 2188 8072 2194 8084
rect 2685 8075 2743 8081
rect 2685 8072 2697 8075
rect 2188 8044 2697 8072
rect 2188 8032 2194 8044
rect 2685 8041 2697 8044
rect 2731 8041 2743 8075
rect 2685 8035 2743 8041
rect 4614 8032 4620 8084
rect 4672 8072 4678 8084
rect 5997 8075 6055 8081
rect 5997 8072 6009 8075
rect 4672 8044 6009 8072
rect 4672 8032 4678 8044
rect 5997 8041 6009 8044
rect 6043 8041 6055 8075
rect 5997 8035 6055 8041
rect 9306 8032 9312 8084
rect 9364 8072 9370 8084
rect 9401 8075 9459 8081
rect 9401 8072 9413 8075
rect 9364 8044 9413 8072
rect 9364 8032 9370 8044
rect 9401 8041 9413 8044
rect 9447 8041 9459 8075
rect 9401 8035 9459 8041
rect 2958 7964 2964 8016
rect 3016 8004 3022 8016
rect 3234 8004 3240 8016
rect 3016 7976 3240 8004
rect 3016 7964 3022 7976
rect 3234 7964 3240 7976
rect 3292 7964 3298 8016
rect 5721 8007 5779 8013
rect 5721 8004 5733 8007
rect 4264 7976 5733 8004
rect 1964 7908 2728 7936
rect 1964 7877 1992 7908
rect 1949 7871 2007 7877
rect 1949 7837 1961 7871
rect 1995 7837 2007 7871
rect 1949 7831 2007 7837
rect 2041 7871 2099 7877
rect 2041 7837 2053 7871
rect 2087 7837 2099 7871
rect 2041 7831 2099 7837
rect 1305 7803 1363 7809
rect 1305 7769 1317 7803
rect 1351 7800 1363 7803
rect 2056 7800 2084 7831
rect 1351 7772 2084 7800
rect 2700 7800 2728 7908
rect 2777 7871 2835 7877
rect 2777 7837 2789 7871
rect 2823 7868 2835 7871
rect 2958 7868 2964 7880
rect 2823 7840 2964 7868
rect 2823 7837 2835 7840
rect 2777 7831 2835 7837
rect 2958 7828 2964 7840
rect 3016 7828 3022 7880
rect 4264 7877 4292 7976
rect 5721 7973 5733 7976
rect 5767 7973 5779 8007
rect 5721 7967 5779 7973
rect 7926 7964 7932 8016
rect 7984 8004 7990 8016
rect 8570 8004 8576 8016
rect 7984 7976 8576 8004
rect 7984 7964 7990 7976
rect 8570 7964 8576 7976
rect 8628 7964 8634 8016
rect 5626 7896 5632 7948
rect 5684 7936 5690 7948
rect 6089 7939 6147 7945
rect 6089 7936 6101 7939
rect 5684 7908 6101 7936
rect 5684 7896 5690 7908
rect 6089 7905 6101 7908
rect 6135 7936 6147 7939
rect 6362 7936 6368 7948
rect 6135 7908 6368 7936
rect 6135 7905 6147 7908
rect 6089 7899 6147 7905
rect 6362 7896 6368 7908
rect 6420 7896 6426 7948
rect 7098 7896 7104 7948
rect 7156 7936 7162 7948
rect 7156 7908 8248 7936
rect 7156 7896 7162 7908
rect 4249 7871 4307 7877
rect 4249 7837 4261 7871
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4341 7871 4399 7877
rect 4341 7837 4353 7871
rect 4387 7837 4399 7871
rect 4341 7831 4399 7837
rect 3421 7803 3479 7809
rect 3421 7800 3433 7803
rect 2700 7772 3433 7800
rect 1351 7769 1363 7772
rect 1305 7763 1363 7769
rect 3421 7769 3433 7772
rect 3467 7769 3479 7803
rect 3421 7763 3479 7769
rect 3605 7803 3663 7809
rect 3605 7769 3617 7803
rect 3651 7800 3663 7803
rect 4356 7800 4384 7831
rect 4430 7828 4436 7880
rect 4488 7868 4494 7880
rect 5077 7871 5135 7877
rect 5077 7868 5089 7871
rect 4488 7840 5089 7868
rect 4488 7828 4494 7840
rect 5077 7837 5089 7840
rect 5123 7837 5135 7871
rect 5077 7831 5135 7837
rect 5718 7828 5724 7880
rect 5776 7868 5782 7880
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5776 7840 5825 7868
rect 5776 7828 5782 7840
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 7466 7828 7472 7880
rect 7524 7828 7530 7880
rect 8220 7877 8248 7908
rect 8205 7871 8263 7877
rect 8205 7837 8217 7871
rect 8251 7837 8263 7871
rect 8205 7831 8263 7837
rect 8573 7871 8631 7877
rect 8573 7837 8585 7871
rect 8619 7868 8631 7871
rect 8662 7868 8668 7880
rect 8619 7840 8668 7868
rect 8619 7837 8631 7840
rect 8573 7831 8631 7837
rect 8662 7828 8668 7840
rect 8720 7828 8726 7880
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 8812 7840 8857 7868
rect 8812 7828 8818 7840
rect 3651 7772 4384 7800
rect 6365 7803 6423 7809
rect 3651 7769 3663 7772
rect 3605 7763 3663 7769
rect 6365 7769 6377 7803
rect 6411 7800 6423 7803
rect 6454 7800 6460 7812
rect 6411 7772 6460 7800
rect 6411 7769 6423 7772
rect 6365 7763 6423 7769
rect 6454 7760 6460 7772
rect 6512 7760 6518 7812
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 4985 7735 5043 7741
rect 4985 7732 4997 7735
rect 3936 7704 4997 7732
rect 3936 7692 3942 7704
rect 4985 7701 4997 7704
rect 5031 7701 5043 7735
rect 4985 7695 5043 7701
rect 7190 7692 7196 7744
rect 7248 7732 7254 7744
rect 7484 7732 7512 7828
rect 7248 7704 7512 7732
rect 7837 7735 7895 7741
rect 7248 7692 7254 7704
rect 7837 7701 7849 7735
rect 7883 7732 7895 7735
rect 7926 7732 7932 7744
rect 7883 7704 7932 7732
rect 7883 7701 7895 7704
rect 7837 7695 7895 7701
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 8110 7732 8116 7744
rect 8071 7704 8116 7732
rect 8110 7692 8116 7704
rect 8168 7692 8174 7744
rect 8294 7732 8300 7744
rect 8255 7704 8300 7732
rect 8294 7692 8300 7704
rect 8352 7692 8358 7744
rect 8386 7692 8392 7744
rect 8444 7732 8450 7744
rect 8444 7704 8489 7732
rect 8444 7692 8450 7704
rect 920 7642 9844 7664
rect 920 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 5194 7642
rect 5246 7590 5258 7642
rect 5310 7590 5322 7642
rect 5374 7590 9844 7642
rect 920 7568 9844 7590
rect 1305 7531 1363 7537
rect 1305 7497 1317 7531
rect 1351 7528 1363 7531
rect 1394 7528 1400 7540
rect 1351 7500 1400 7528
rect 1351 7497 1363 7500
rect 1305 7491 1363 7497
rect 1394 7488 1400 7500
rect 1452 7488 1458 7540
rect 3418 7488 3424 7540
rect 3476 7528 3482 7540
rect 5626 7528 5632 7540
rect 3476 7500 5632 7528
rect 3476 7488 3482 7500
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 5917 7531 5975 7537
rect 5917 7497 5929 7531
rect 5963 7528 5975 7531
rect 8386 7528 8392 7540
rect 5963 7500 8392 7528
rect 5963 7497 5975 7500
rect 5917 7491 5975 7497
rect 8386 7488 8392 7500
rect 8444 7488 8450 7540
rect 1412 7460 1440 7488
rect 1412 7446 1978 7460
rect 1412 7432 1992 7446
rect 1964 7324 1992 7432
rect 3142 7420 3148 7472
rect 3200 7460 3206 7472
rect 5442 7460 5448 7472
rect 3200 7432 3556 7460
rect 5014 7432 5448 7460
rect 3200 7420 3206 7432
rect 3528 7401 3556 7432
rect 5442 7420 5448 7432
rect 5500 7420 5506 7472
rect 7466 7420 7472 7472
rect 7524 7420 7530 7472
rect 3513 7395 3571 7401
rect 3513 7361 3525 7395
rect 3559 7361 3571 7395
rect 3878 7392 3884 7404
rect 3839 7364 3884 7392
rect 3513 7355 3571 7361
rect 3878 7352 3884 7364
rect 3936 7352 3942 7404
rect 4798 7352 4804 7404
rect 4856 7392 4862 7404
rect 5353 7395 5411 7401
rect 5353 7392 5365 7395
rect 4856 7364 5365 7392
rect 4856 7352 4862 7364
rect 5353 7361 5365 7364
rect 5399 7361 5411 7395
rect 5353 7355 5411 7361
rect 6365 7395 6423 7401
rect 6365 7361 6377 7395
rect 6411 7392 6423 7395
rect 6822 7392 6828 7404
rect 6411 7364 6828 7392
rect 6411 7361 6423 7364
rect 6365 7355 6423 7361
rect 6822 7352 6828 7364
rect 6880 7352 6886 7404
rect 8202 7392 8208 7404
rect 8163 7364 8208 7392
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 8404 7392 8432 7488
rect 8941 7395 8999 7401
rect 8941 7392 8953 7395
rect 8404 7364 8953 7392
rect 8941 7361 8953 7364
rect 8987 7361 8999 7395
rect 8941 7355 8999 7361
rect 2406 7324 2412 7336
rect 1964 7296 2412 7324
rect 2406 7284 2412 7296
rect 2464 7284 2470 7336
rect 3050 7284 3056 7336
rect 3108 7324 3114 7336
rect 3145 7327 3203 7333
rect 3145 7324 3157 7327
rect 3108 7296 3157 7324
rect 3108 7284 3114 7296
rect 3145 7293 3157 7296
rect 3191 7293 3203 7327
rect 3418 7324 3424 7336
rect 3379 7296 3424 7324
rect 3145 7287 3203 7293
rect 3418 7284 3424 7296
rect 3476 7284 3482 7336
rect 6733 7327 6791 7333
rect 6733 7293 6745 7327
rect 6779 7324 6791 7327
rect 7006 7324 7012 7336
rect 6779 7296 7012 7324
rect 6779 7293 6791 7296
rect 6733 7287 6791 7293
rect 7006 7284 7012 7296
rect 7064 7284 7070 7336
rect 4798 7216 4804 7268
rect 4856 7256 4862 7268
rect 4982 7256 4988 7268
rect 4856 7228 4988 7256
rect 4856 7216 4862 7228
rect 4982 7216 4988 7228
rect 5040 7256 5046 7268
rect 6181 7259 6239 7265
rect 6181 7256 6193 7259
rect 5040 7228 6193 7256
rect 5040 7216 5046 7228
rect 6181 7225 6193 7228
rect 6227 7225 6239 7259
rect 6181 7219 6239 7225
rect 1670 7188 1676 7200
rect 1631 7160 1676 7188
rect 1670 7148 1676 7160
rect 1728 7148 1734 7200
rect 8294 7148 8300 7200
rect 8352 7188 8358 7200
rect 8389 7191 8447 7197
rect 8389 7188 8401 7191
rect 8352 7160 8401 7188
rect 8352 7148 8358 7160
rect 8389 7157 8401 7160
rect 8435 7157 8447 7191
rect 8389 7151 8447 7157
rect 8769 7191 8827 7197
rect 8769 7157 8781 7191
rect 8815 7188 8827 7191
rect 8938 7188 8944 7200
rect 8815 7160 8944 7188
rect 8815 7157 8827 7160
rect 8769 7151 8827 7157
rect 8938 7148 8944 7160
rect 8996 7148 9002 7200
rect 9030 7148 9036 7200
rect 9088 7188 9094 7200
rect 9088 7160 9133 7188
rect 9088 7148 9094 7160
rect 9306 7148 9312 7200
rect 9364 7188 9370 7200
rect 9401 7191 9459 7197
rect 9401 7188 9413 7191
rect 9364 7160 9413 7188
rect 9364 7148 9370 7160
rect 9401 7157 9413 7160
rect 9447 7157 9459 7191
rect 9401 7151 9459 7157
rect 920 7098 9844 7120
rect 920 7046 2566 7098
rect 2618 7046 2630 7098
rect 2682 7046 2694 7098
rect 2746 7046 2758 7098
rect 2810 7046 2822 7098
rect 2874 7046 7566 7098
rect 7618 7046 7630 7098
rect 7682 7046 7694 7098
rect 7746 7046 7758 7098
rect 7810 7046 7822 7098
rect 7874 7046 9844 7098
rect 920 7024 9844 7046
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 2795 6987 2853 6993
rect 2795 6984 2807 6987
rect 1728 6956 2807 6984
rect 1728 6944 1734 6956
rect 2795 6953 2807 6956
rect 2841 6984 2853 6987
rect 4430 6984 4436 6996
rect 2841 6956 4436 6984
rect 2841 6953 2853 6956
rect 2795 6947 2853 6953
rect 4430 6944 4436 6956
rect 4488 6944 4494 6996
rect 4154 6916 4160 6928
rect 4080 6888 4160 6916
rect 3053 6851 3111 6857
rect 3053 6817 3065 6851
rect 3099 6848 3111 6851
rect 3418 6848 3424 6860
rect 3099 6820 3424 6848
rect 3099 6817 3111 6820
rect 3053 6811 3111 6817
rect 3418 6808 3424 6820
rect 3476 6808 3482 6860
rect 3237 6783 3295 6789
rect 3237 6749 3249 6783
rect 3283 6780 3295 6783
rect 4080 6780 4108 6888
rect 4154 6876 4160 6888
rect 4212 6876 4218 6928
rect 5721 6919 5779 6925
rect 5721 6916 5733 6919
rect 4264 6888 5733 6916
rect 4264 6789 4292 6888
rect 5721 6885 5733 6888
rect 5767 6885 5779 6919
rect 5721 6879 5779 6885
rect 7190 6876 7196 6928
rect 7248 6916 7254 6928
rect 8110 6916 8116 6928
rect 7248 6888 8116 6916
rect 7248 6876 7254 6888
rect 8110 6876 8116 6888
rect 8168 6876 8174 6928
rect 6270 6848 6276 6860
rect 6231 6820 6276 6848
rect 6270 6808 6276 6820
rect 6328 6808 6334 6860
rect 7926 6808 7932 6860
rect 7984 6848 7990 6860
rect 7984 6820 8616 6848
rect 7984 6808 7990 6820
rect 3283 6752 4108 6780
rect 4249 6783 4307 6789
rect 3283 6749 3295 6752
rect 3237 6743 3295 6749
rect 4249 6749 4261 6783
rect 4295 6749 4307 6783
rect 4249 6743 4307 6749
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6749 4399 6783
rect 4341 6743 4399 6749
rect 2498 6712 2504 6724
rect 2346 6684 2504 6712
rect 2498 6672 2504 6684
rect 2556 6712 2562 6724
rect 2682 6712 2688 6724
rect 2556 6684 2688 6712
rect 2556 6672 2562 6684
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 3605 6715 3663 6721
rect 3605 6681 3617 6715
rect 3651 6712 3663 6715
rect 4356 6712 4384 6743
rect 5074 6740 5080 6792
rect 5132 6780 5138 6792
rect 5132 6752 5177 6780
rect 5132 6740 5138 6752
rect 5810 6740 5816 6792
rect 5868 6780 5874 6792
rect 5997 6783 6055 6789
rect 5997 6780 6009 6783
rect 5868 6752 6009 6780
rect 5868 6740 5874 6752
rect 5997 6749 6009 6752
rect 6043 6749 6055 6783
rect 5997 6743 6055 6749
rect 7837 6783 7895 6789
rect 7837 6749 7849 6783
rect 7883 6780 7895 6783
rect 8018 6780 8024 6792
rect 7883 6752 8024 6780
rect 7883 6749 7895 6752
rect 7837 6743 7895 6749
rect 8018 6740 8024 6752
rect 8076 6740 8082 6792
rect 8588 6789 8616 6820
rect 8573 6783 8631 6789
rect 8573 6749 8585 6783
rect 8619 6749 8631 6783
rect 8573 6743 8631 6749
rect 9122 6740 9128 6792
rect 9180 6780 9186 6792
rect 9493 6783 9551 6789
rect 9493 6780 9505 6783
rect 9180 6752 9505 6780
rect 9180 6740 9186 6752
rect 9493 6749 9505 6752
rect 9539 6749 9551 6783
rect 9493 6743 9551 6749
rect 3651 6684 4384 6712
rect 3651 6681 3663 6684
rect 3605 6675 3663 6681
rect 7190 6672 7196 6724
rect 7248 6712 7254 6724
rect 8849 6715 8907 6721
rect 8849 6712 8861 6715
rect 7248 6684 8861 6712
rect 7248 6672 7254 6684
rect 8849 6681 8861 6684
rect 8895 6681 8907 6715
rect 8849 6675 8907 6681
rect 1305 6647 1363 6653
rect 1305 6613 1317 6647
rect 1351 6644 1363 6647
rect 1486 6644 1492 6656
rect 1351 6616 1492 6644
rect 1351 6613 1363 6616
rect 1305 6607 1363 6613
rect 1486 6604 1492 6616
rect 1544 6644 1550 6656
rect 2958 6644 2964 6656
rect 1544 6616 2964 6644
rect 1544 6604 1550 6616
rect 2958 6604 2964 6616
rect 3016 6604 3022 6656
rect 3418 6644 3424 6656
rect 3379 6616 3424 6644
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 4062 6604 4068 6656
rect 4120 6644 4126 6656
rect 4985 6647 5043 6653
rect 4985 6644 4997 6647
rect 4120 6616 4997 6644
rect 4120 6604 4126 6616
rect 4985 6613 4997 6616
rect 5031 6613 5043 6647
rect 4985 6607 5043 6613
rect 5810 6604 5816 6656
rect 5868 6644 5874 6656
rect 5868 6616 5913 6644
rect 5868 6604 5874 6616
rect 6362 6604 6368 6656
rect 6420 6644 6426 6656
rect 6822 6644 6828 6656
rect 6420 6616 6828 6644
rect 6420 6604 6426 6616
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7098 6604 7104 6656
rect 7156 6644 7162 6656
rect 7929 6647 7987 6653
rect 7929 6644 7941 6647
rect 7156 6616 7941 6644
rect 7156 6604 7162 6616
rect 7929 6613 7941 6616
rect 7975 6613 7987 6647
rect 7929 6607 7987 6613
rect 920 6554 9844 6576
rect 920 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 5194 6554
rect 5246 6502 5258 6554
rect 5310 6502 5322 6554
rect 5374 6502 9844 6554
rect 920 6480 9844 6502
rect 5905 6443 5963 6449
rect 5905 6440 5917 6443
rect 3252 6412 5917 6440
rect 1486 6332 1492 6384
rect 1544 6372 1550 6384
rect 1581 6375 1639 6381
rect 1581 6372 1593 6375
rect 1544 6344 1593 6372
rect 1544 6332 1550 6344
rect 1581 6341 1593 6344
rect 1627 6341 1639 6375
rect 1581 6335 1639 6341
rect 2682 6264 2688 6316
rect 2740 6304 2746 6316
rect 3142 6304 3148 6316
rect 2740 6276 3148 6304
rect 2740 6264 2746 6276
rect 3142 6264 3148 6276
rect 3200 6264 3206 6316
rect 3252 6313 3280 6412
rect 5905 6409 5917 6412
rect 5951 6409 5963 6443
rect 7006 6440 7012 6452
rect 5905 6403 5963 6409
rect 6564 6412 7012 6440
rect 3970 6332 3976 6384
rect 4028 6332 4034 6384
rect 3237 6307 3295 6313
rect 3237 6273 3249 6307
rect 3283 6273 3295 6307
rect 3237 6267 3295 6273
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5810 6304 5816 6316
rect 5123 6276 5816 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 5810 6264 5816 6276
rect 5868 6264 5874 6316
rect 5994 6304 6000 6316
rect 5955 6276 6000 6304
rect 5994 6264 6000 6276
rect 6052 6264 6058 6316
rect 6178 6264 6184 6316
rect 6236 6304 6242 6316
rect 6564 6313 6592 6412
rect 7006 6400 7012 6412
rect 7064 6440 7070 6452
rect 7834 6440 7840 6452
rect 7064 6412 7840 6440
rect 7064 6400 7070 6412
rect 7834 6400 7840 6412
rect 7892 6400 7898 6452
rect 6822 6332 6828 6384
rect 6880 6372 6886 6384
rect 7653 6375 7711 6381
rect 6880 6344 7420 6372
rect 6880 6332 6886 6344
rect 6365 6307 6423 6313
rect 6365 6304 6377 6307
rect 6236 6276 6377 6304
rect 6236 6264 6242 6276
rect 6365 6273 6377 6276
rect 6411 6273 6423 6307
rect 6365 6267 6423 6273
rect 6549 6307 6607 6313
rect 6549 6273 6561 6307
rect 6595 6273 6607 6307
rect 6549 6267 6607 6273
rect 6733 6307 6791 6313
rect 6733 6273 6745 6307
rect 6779 6273 6791 6307
rect 7006 6304 7012 6316
rect 6967 6276 7012 6304
rect 6733 6267 6791 6273
rect 1302 6236 1308 6248
rect 1263 6208 1308 6236
rect 1302 6196 1308 6208
rect 1360 6196 1366 6248
rect 3602 6236 3608 6248
rect 3563 6208 3608 6236
rect 3602 6196 3608 6208
rect 3660 6196 3666 6248
rect 5442 6128 5448 6180
rect 5500 6168 5506 6180
rect 6181 6171 6239 6177
rect 6181 6168 6193 6171
rect 5500 6140 6193 6168
rect 5500 6128 5506 6140
rect 6181 6137 6193 6140
rect 6227 6137 6239 6171
rect 6748 6168 6776 6267
rect 7006 6264 7012 6276
rect 7064 6264 7070 6316
rect 7392 6313 7420 6344
rect 7653 6341 7665 6375
rect 7699 6372 7711 6375
rect 7926 6372 7932 6384
rect 7699 6344 7932 6372
rect 7699 6341 7711 6344
rect 7653 6335 7711 6341
rect 7926 6332 7932 6344
rect 7984 6332 7990 6384
rect 8110 6332 8116 6384
rect 8168 6332 8174 6384
rect 7285 6307 7343 6313
rect 7285 6273 7297 6307
rect 7331 6273 7343 6307
rect 7285 6267 7343 6273
rect 7377 6307 7435 6313
rect 7377 6273 7389 6307
rect 7423 6273 7435 6307
rect 7377 6267 7435 6273
rect 6914 6236 6920 6248
rect 6875 6208 6920 6236
rect 6914 6196 6920 6208
rect 6972 6196 6978 6248
rect 7300 6236 7328 6267
rect 9398 6264 9404 6316
rect 9456 6304 9462 6316
rect 9493 6307 9551 6313
rect 9493 6304 9505 6307
rect 9456 6276 9505 6304
rect 9456 6264 9462 6276
rect 9493 6273 9505 6276
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 8110 6236 8116 6248
rect 7300 6208 8116 6236
rect 8110 6196 8116 6208
rect 8168 6196 8174 6248
rect 8202 6196 8208 6248
rect 8260 6236 8266 6248
rect 8260 6208 9352 6236
rect 8260 6196 8266 6208
rect 7282 6168 7288 6180
rect 6748 6140 7288 6168
rect 6181 6131 6239 6137
rect 7282 6128 7288 6140
rect 7340 6128 7346 6180
rect 9324 6177 9352 6208
rect 9309 6171 9367 6177
rect 9309 6137 9321 6171
rect 9355 6137 9367 6171
rect 9309 6131 9367 6137
rect 1946 6060 1952 6112
rect 2004 6100 2010 6112
rect 3053 6103 3111 6109
rect 3053 6100 3065 6103
rect 2004 6072 3065 6100
rect 2004 6060 2010 6072
rect 3053 6069 3065 6072
rect 3099 6100 3111 6103
rect 4982 6100 4988 6112
rect 3099 6072 4988 6100
rect 3099 6069 3111 6072
rect 3053 6063 3111 6069
rect 4982 6060 4988 6072
rect 5040 6060 5046 6112
rect 5641 6103 5699 6109
rect 5641 6069 5653 6103
rect 5687 6100 5699 6103
rect 6822 6100 6828 6112
rect 5687 6072 6828 6100
rect 5687 6069 5699 6072
rect 5641 6063 5699 6069
rect 6822 6060 6828 6072
rect 6880 6060 6886 6112
rect 9122 6100 9128 6112
rect 9083 6072 9128 6100
rect 9122 6060 9128 6072
rect 9180 6060 9186 6112
rect 920 6010 9844 6032
rect 920 5958 2566 6010
rect 2618 5958 2630 6010
rect 2682 5958 2694 6010
rect 2746 5958 2758 6010
rect 2810 5958 2822 6010
rect 2874 5958 7566 6010
rect 7618 5958 7630 6010
rect 7682 5958 7694 6010
rect 7746 5958 7758 6010
rect 7810 5958 7822 6010
rect 7874 5958 9844 6010
rect 920 5936 9844 5958
rect 3697 5899 3755 5905
rect 3697 5896 3709 5899
rect 1228 5868 3709 5896
rect 1228 5692 1256 5868
rect 3697 5865 3709 5868
rect 3743 5865 3755 5899
rect 3697 5859 3755 5865
rect 4065 5899 4123 5905
rect 4065 5865 4077 5899
rect 4111 5865 4123 5899
rect 4065 5859 4123 5865
rect 1302 5788 1308 5840
rect 1360 5788 1366 5840
rect 4080 5828 4108 5859
rect 4338 5856 4344 5908
rect 4396 5896 4402 5908
rect 5442 5896 5448 5908
rect 4396 5868 5448 5896
rect 4396 5856 4402 5868
rect 5442 5856 5448 5868
rect 5500 5896 5506 5908
rect 5537 5899 5595 5905
rect 5537 5896 5549 5899
rect 5500 5868 5549 5896
rect 5500 5856 5506 5868
rect 5537 5865 5549 5868
rect 5583 5865 5595 5899
rect 5537 5859 5595 5865
rect 6273 5899 6331 5905
rect 6273 5865 6285 5899
rect 6319 5896 6331 5899
rect 6914 5896 6920 5908
rect 6319 5868 6920 5896
rect 6319 5865 6331 5868
rect 6273 5859 6331 5865
rect 4614 5828 4620 5840
rect 4080 5800 4620 5828
rect 4614 5788 4620 5800
rect 4672 5828 4678 5840
rect 6288 5828 6316 5859
rect 6914 5856 6920 5868
rect 6972 5856 6978 5908
rect 7006 5856 7012 5908
rect 7064 5896 7070 5908
rect 7745 5899 7803 5905
rect 7745 5896 7757 5899
rect 7064 5868 7757 5896
rect 7064 5856 7070 5868
rect 7745 5865 7757 5868
rect 7791 5865 7803 5899
rect 7745 5859 7803 5865
rect 8110 5856 8116 5908
rect 8168 5896 8174 5908
rect 8849 5899 8907 5905
rect 8849 5896 8861 5899
rect 8168 5868 8861 5896
rect 8168 5856 8174 5868
rect 8849 5865 8861 5868
rect 8895 5865 8907 5899
rect 8849 5859 8907 5865
rect 8938 5856 8944 5908
rect 8996 5896 9002 5908
rect 11514 5896 11520 5908
rect 8996 5868 11520 5896
rect 8996 5856 9002 5868
rect 11514 5856 11520 5868
rect 11572 5856 11578 5908
rect 4672 5800 6316 5828
rect 6641 5831 6699 5837
rect 4672 5788 4678 5800
rect 6641 5797 6653 5831
rect 6687 5828 6699 5831
rect 9490 5828 9496 5840
rect 6687 5800 9496 5828
rect 6687 5797 6699 5800
rect 6641 5791 6699 5797
rect 9490 5788 9496 5800
rect 9548 5788 9554 5840
rect 1320 5760 1348 5788
rect 1581 5763 1639 5769
rect 1581 5760 1593 5763
rect 1320 5732 1593 5760
rect 1581 5729 1593 5732
rect 1627 5760 1639 5763
rect 1627 5732 3372 5760
rect 1627 5729 1639 5732
rect 1581 5723 1639 5729
rect 1305 5695 1363 5701
rect 1305 5692 1317 5695
rect 1228 5664 1317 5692
rect 1305 5661 1317 5664
rect 1351 5661 1363 5695
rect 3344 5692 3372 5732
rect 3418 5720 3424 5772
rect 3476 5760 3482 5772
rect 6730 5760 6736 5772
rect 3476 5732 4292 5760
rect 3476 5720 3482 5732
rect 3878 5692 3884 5704
rect 3344 5664 3884 5692
rect 1305 5655 1363 5661
rect 3878 5652 3884 5664
rect 3936 5652 3942 5704
rect 4264 5701 4292 5732
rect 6196 5732 6736 5760
rect 6196 5701 6224 5732
rect 6730 5720 6736 5732
rect 6788 5720 6794 5772
rect 7285 5763 7343 5769
rect 7285 5729 7297 5763
rect 7331 5760 7343 5763
rect 8846 5760 8852 5772
rect 7331 5732 8064 5760
rect 7331 5729 7343 5732
rect 7285 5723 7343 5729
rect 4157 5695 4215 5701
rect 4157 5661 4169 5695
rect 4203 5661 4215 5695
rect 4157 5655 4215 5661
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 6181 5695 6239 5701
rect 6181 5661 6193 5695
rect 6227 5661 6239 5695
rect 6181 5655 6239 5661
rect 1857 5627 1915 5633
rect 1857 5593 1869 5627
rect 1903 5624 1915 5627
rect 1946 5624 1952 5636
rect 1903 5596 1952 5624
rect 1903 5593 1915 5596
rect 1857 5587 1915 5593
rect 1946 5584 1952 5596
rect 2004 5584 2010 5636
rect 3142 5624 3148 5636
rect 3082 5596 3148 5624
rect 3142 5584 3148 5596
rect 3200 5584 3206 5636
rect 3970 5624 3976 5636
rect 3252 5596 3976 5624
rect 1489 5559 1547 5565
rect 1489 5525 1501 5559
rect 1535 5556 1547 5559
rect 3252 5556 3280 5596
rect 3970 5584 3976 5596
rect 4028 5584 4034 5636
rect 4172 5624 4200 5655
rect 6546 5652 6552 5704
rect 6604 5692 6610 5704
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 6604 5664 6837 5692
rect 6604 5652 6610 5664
rect 6825 5661 6837 5664
rect 6871 5661 6883 5695
rect 6825 5655 6883 5661
rect 7469 5695 7527 5701
rect 7469 5661 7481 5695
rect 7515 5661 7527 5695
rect 7469 5655 7527 5661
rect 7745 5695 7803 5701
rect 7745 5661 7757 5695
rect 7791 5692 7803 5695
rect 7926 5692 7932 5704
rect 7791 5664 7932 5692
rect 7791 5661 7803 5664
rect 7745 5655 7803 5661
rect 4798 5624 4804 5636
rect 4172 5596 4804 5624
rect 4798 5584 4804 5596
rect 4856 5584 4862 5636
rect 5718 5584 5724 5636
rect 5776 5624 5782 5636
rect 6086 5624 6092 5636
rect 5776 5596 6092 5624
rect 5776 5584 5782 5596
rect 6086 5584 6092 5596
rect 6144 5624 6150 5636
rect 7484 5624 7512 5655
rect 7926 5652 7932 5664
rect 7984 5652 7990 5704
rect 6144 5596 7512 5624
rect 8036 5624 8064 5732
rect 8128 5732 8852 5760
rect 8128 5701 8156 5732
rect 8846 5720 8852 5732
rect 8904 5760 8910 5772
rect 9217 5763 9275 5769
rect 9217 5760 9229 5763
rect 8904 5732 9229 5760
rect 8904 5720 8910 5732
rect 9217 5729 9229 5732
rect 9263 5729 9275 5763
rect 9217 5723 9275 5729
rect 8113 5695 8171 5701
rect 8113 5661 8125 5695
rect 8159 5661 8171 5695
rect 8294 5692 8300 5704
rect 8255 5664 8300 5692
rect 8113 5655 8171 5661
rect 8294 5652 8300 5664
rect 8352 5652 8358 5704
rect 8573 5695 8631 5701
rect 8573 5661 8585 5695
rect 8619 5661 8631 5695
rect 9030 5692 9036 5704
rect 8991 5664 9036 5692
rect 8573 5655 8631 5661
rect 8202 5624 8208 5636
rect 8036 5596 8208 5624
rect 6144 5584 6150 5596
rect 8202 5584 8208 5596
rect 8260 5584 8266 5636
rect 8588 5624 8616 5655
rect 9030 5652 9036 5664
rect 9088 5652 9094 5704
rect 9309 5695 9367 5701
rect 9309 5661 9321 5695
rect 9355 5661 9367 5695
rect 9309 5655 9367 5661
rect 8754 5624 8760 5636
rect 8588 5596 8760 5624
rect 8754 5584 8760 5596
rect 8812 5624 8818 5636
rect 9324 5624 9352 5655
rect 8812 5596 9352 5624
rect 8812 5584 8818 5596
rect 1535 5528 3280 5556
rect 1535 5525 1547 5528
rect 1489 5519 1547 5525
rect 3326 5516 3332 5568
rect 3384 5556 3390 5568
rect 3384 5528 3429 5556
rect 3384 5516 3390 5528
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 7282 5556 7288 5568
rect 6604 5528 7288 5556
rect 6604 5516 6610 5528
rect 7282 5516 7288 5528
rect 7340 5516 7346 5568
rect 7653 5559 7711 5565
rect 7653 5525 7665 5559
rect 7699 5556 7711 5559
rect 7926 5556 7932 5568
rect 7699 5528 7932 5556
rect 7699 5525 7711 5528
rect 7653 5519 7711 5525
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 8294 5516 8300 5568
rect 8352 5556 8358 5568
rect 8570 5556 8576 5568
rect 8352 5528 8576 5556
rect 8352 5516 8358 5528
rect 8570 5516 8576 5528
rect 8628 5516 8634 5568
rect 9214 5516 9220 5568
rect 9272 5556 9278 5568
rect 9401 5559 9459 5565
rect 9401 5556 9413 5559
rect 9272 5528 9413 5556
rect 9272 5516 9278 5528
rect 9401 5525 9413 5528
rect 9447 5525 9459 5559
rect 9401 5519 9459 5525
rect 920 5466 9844 5488
rect 920 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 5194 5466
rect 5246 5414 5258 5466
rect 5310 5414 5322 5466
rect 5374 5414 9844 5466
rect 920 5392 9844 5414
rect 3602 5312 3608 5364
rect 3660 5352 3666 5364
rect 4801 5355 4859 5361
rect 4801 5352 4813 5355
rect 3660 5324 4813 5352
rect 3660 5312 3666 5324
rect 4801 5321 4813 5324
rect 4847 5321 4859 5355
rect 5718 5352 5724 5364
rect 5631 5324 5724 5352
rect 4801 5315 4859 5321
rect 5718 5312 5724 5324
rect 5776 5352 5782 5364
rect 5902 5352 5908 5364
rect 5776 5324 5908 5352
rect 5776 5312 5782 5324
rect 5902 5312 5908 5324
rect 5960 5312 5966 5364
rect 6730 5312 6736 5364
rect 6788 5352 6794 5364
rect 6788 5324 7512 5352
rect 6788 5312 6794 5324
rect 5077 5287 5135 5293
rect 5077 5253 5089 5287
rect 5123 5284 5135 5287
rect 6270 5284 6276 5296
rect 5123 5256 6276 5284
rect 5123 5253 5135 5256
rect 5077 5247 5135 5253
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 7009 5287 7067 5293
rect 7009 5253 7021 5287
rect 7055 5284 7067 5287
rect 7374 5284 7380 5296
rect 7055 5256 7380 5284
rect 7055 5253 7067 5256
rect 7009 5247 7067 5253
rect 7374 5244 7380 5256
rect 7432 5244 7438 5296
rect 7484 5284 7512 5324
rect 7650 5312 7656 5364
rect 7708 5352 7714 5364
rect 9309 5355 9367 5361
rect 9309 5352 9321 5355
rect 7708 5324 9321 5352
rect 7708 5312 7714 5324
rect 9309 5321 9321 5324
rect 9355 5321 9367 5355
rect 9309 5315 9367 5321
rect 7745 5287 7803 5293
rect 7745 5284 7757 5287
rect 7484 5256 7757 5284
rect 7745 5253 7757 5256
rect 7791 5253 7803 5287
rect 8481 5287 8539 5293
rect 8481 5284 8493 5287
rect 7745 5247 7803 5253
rect 7944 5256 8493 5284
rect 7944 5228 7972 5256
rect 8481 5253 8493 5256
rect 8527 5253 8539 5287
rect 8846 5284 8852 5296
rect 8807 5256 8852 5284
rect 8481 5247 8539 5253
rect 8846 5244 8852 5256
rect 8904 5244 8910 5296
rect 3418 5216 3424 5228
rect 3379 5188 3424 5216
rect 3418 5176 3424 5188
rect 3476 5176 3482 5228
rect 4065 5219 4123 5225
rect 4065 5185 4077 5219
rect 4111 5216 4123 5219
rect 4157 5219 4215 5225
rect 4157 5216 4169 5219
rect 4111 5188 4169 5216
rect 4111 5185 4123 5188
rect 4065 5179 4123 5185
rect 4157 5185 4169 5188
rect 4203 5185 4215 5219
rect 4157 5179 4215 5185
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 7101 5219 7159 5225
rect 7101 5216 7113 5219
rect 6696 5188 7113 5216
rect 6696 5176 6702 5188
rect 7101 5185 7113 5188
rect 7147 5185 7159 5219
rect 7926 5216 7932 5228
rect 7887 5188 7932 5216
rect 7101 5179 7159 5185
rect 7926 5176 7932 5188
rect 7984 5176 7990 5228
rect 8297 5219 8355 5225
rect 8297 5216 8309 5219
rect 8036 5188 8309 5216
rect 7282 5108 7288 5160
rect 7340 5148 7346 5160
rect 8036 5148 8064 5188
rect 8297 5185 8309 5188
rect 8343 5185 8355 5219
rect 8297 5179 8355 5185
rect 8386 5176 8392 5228
rect 8444 5216 8450 5228
rect 8570 5216 8576 5228
rect 8444 5188 8576 5216
rect 8444 5176 8450 5188
rect 8570 5176 8576 5188
rect 8628 5216 8634 5228
rect 8941 5219 8999 5225
rect 8941 5216 8953 5219
rect 8628 5188 8953 5216
rect 8628 5176 8634 5188
rect 8941 5185 8953 5188
rect 8987 5185 8999 5219
rect 9214 5216 9220 5228
rect 9175 5188 9220 5216
rect 8941 5179 8999 5185
rect 9214 5176 9220 5188
rect 9272 5176 9278 5228
rect 9490 5216 9496 5228
rect 9451 5188 9496 5216
rect 9490 5176 9496 5188
rect 9548 5176 9554 5228
rect 7340 5120 8064 5148
rect 8113 5151 8171 5157
rect 7340 5108 7346 5120
rect 8113 5117 8125 5151
rect 8159 5148 8171 5151
rect 9398 5148 9404 5160
rect 8159 5120 9404 5148
rect 8159 5117 8171 5120
rect 8113 5111 8171 5117
rect 9398 5108 9404 5120
rect 9456 5108 9462 5160
rect 4154 5040 4160 5092
rect 4212 5080 4218 5092
rect 4893 5083 4951 5089
rect 4893 5080 4905 5083
rect 4212 5052 4905 5080
rect 4212 5040 4218 5052
rect 4893 5049 4905 5052
rect 4939 5049 4951 5083
rect 4893 5043 4951 5049
rect 8665 5083 8723 5089
rect 8665 5049 8677 5083
rect 8711 5080 8723 5083
rect 8938 5080 8944 5092
rect 8711 5052 8944 5080
rect 8711 5049 8723 5052
rect 8665 5043 8723 5049
rect 8938 5040 8944 5052
rect 8996 5040 9002 5092
rect 3694 4972 3700 5024
rect 3752 5012 3758 5024
rect 4522 5012 4528 5024
rect 3752 4984 4528 5012
rect 3752 4972 3758 4984
rect 4522 4972 4528 4984
rect 4580 5012 4586 5024
rect 5350 5012 5356 5024
rect 4580 4984 5356 5012
rect 4580 4972 4586 4984
rect 5350 4972 5356 4984
rect 5408 5012 5414 5024
rect 5994 5012 6000 5024
rect 5408 4984 6000 5012
rect 5408 4972 5414 4984
rect 5994 4972 6000 4984
rect 6052 4972 6058 5024
rect 6914 4972 6920 5024
rect 6972 5012 6978 5024
rect 7193 5015 7251 5021
rect 7193 5012 7205 5015
rect 6972 4984 7205 5012
rect 6972 4972 6978 4984
rect 7193 4981 7205 4984
rect 7239 4981 7251 5015
rect 7193 4975 7251 4981
rect 7561 5015 7619 5021
rect 7561 4981 7573 5015
rect 7607 5012 7619 5015
rect 7926 5012 7932 5024
rect 7607 4984 7932 5012
rect 7607 4981 7619 4984
rect 7561 4975 7619 4981
rect 7926 4972 7932 4984
rect 7984 4972 7990 5024
rect 3036 4922 9844 4944
rect 3036 4870 7566 4922
rect 7618 4870 7630 4922
rect 7682 4870 7694 4922
rect 7746 4870 7758 4922
rect 7810 4870 7822 4922
rect 7874 4870 9844 4922
rect 3036 4848 9844 4870
rect 3418 4808 3424 4820
rect 3379 4780 3424 4808
rect 3418 4768 3424 4780
rect 3476 4768 3482 4820
rect 4433 4811 4491 4817
rect 4433 4808 4445 4811
rect 3712 4780 4445 4808
rect 3234 4700 3240 4752
rect 3292 4740 3298 4752
rect 3712 4740 3740 4780
rect 4433 4777 4445 4780
rect 4479 4808 4491 4811
rect 5077 4811 5135 4817
rect 5077 4808 5089 4811
rect 4479 4780 5089 4808
rect 4479 4777 4491 4780
rect 4433 4771 4491 4777
rect 5077 4777 5089 4780
rect 5123 4808 5135 4811
rect 5813 4811 5871 4817
rect 5813 4808 5825 4811
rect 5123 4780 5825 4808
rect 5123 4777 5135 4780
rect 5077 4771 5135 4777
rect 5813 4777 5825 4780
rect 5859 4777 5871 4811
rect 5813 4771 5871 4777
rect 8662 4768 8668 4820
rect 8720 4808 8726 4820
rect 9125 4811 9183 4817
rect 9125 4808 9137 4811
rect 8720 4780 9137 4808
rect 8720 4768 8726 4780
rect 9125 4777 9137 4780
rect 9171 4777 9183 4811
rect 9125 4771 9183 4777
rect 3292 4712 3740 4740
rect 3292 4700 3298 4712
rect 4062 4700 4068 4752
rect 4120 4700 4126 4752
rect 4798 4700 4804 4752
rect 4856 4740 4862 4752
rect 5537 4743 5595 4749
rect 5537 4740 5549 4743
rect 4856 4712 5549 4740
rect 4856 4700 4862 4712
rect 5537 4709 5549 4712
rect 5583 4709 5595 4743
rect 5537 4703 5595 4709
rect 4080 4672 4108 4700
rect 6825 4675 6883 4681
rect 4080 4644 5764 4672
rect 3326 4564 3332 4616
rect 3384 4604 3390 4616
rect 3970 4604 3976 4616
rect 3384 4576 3976 4604
rect 3384 4564 3390 4576
rect 3970 4564 3976 4576
rect 4028 4604 4034 4616
rect 4065 4607 4123 4613
rect 4065 4604 4077 4607
rect 4028 4576 4077 4604
rect 4028 4564 4034 4576
rect 4065 4573 4077 4576
rect 4111 4573 4123 4607
rect 4706 4604 4712 4616
rect 4667 4576 4712 4604
rect 4065 4567 4123 4573
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 5350 4604 5356 4616
rect 5311 4576 5356 4604
rect 5350 4564 5356 4576
rect 5408 4564 5414 4616
rect 5736 4613 5764 4644
rect 6825 4641 6837 4675
rect 6871 4672 6883 4675
rect 7098 4672 7104 4684
rect 6871 4644 7104 4672
rect 6871 4641 6883 4644
rect 6825 4635 6883 4641
rect 7098 4632 7104 4644
rect 7156 4632 7162 4684
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 6454 4604 6460 4616
rect 6415 4576 6460 4604
rect 5721 4567 5779 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 8294 4604 8300 4616
rect 8255 4576 8300 4604
rect 8294 4564 8300 4576
rect 8352 4564 8358 4616
rect 9122 4564 9128 4616
rect 9180 4604 9186 4616
rect 9309 4607 9367 4613
rect 9309 4604 9321 4607
rect 9180 4576 9321 4604
rect 9180 4564 9186 4576
rect 9309 4573 9321 4576
rect 9355 4573 9367 4607
rect 9309 4567 9367 4573
rect 9398 4564 9404 4616
rect 9456 4604 9462 4616
rect 9456 4576 9501 4604
rect 9456 4564 9462 4576
rect 4430 4496 4436 4548
rect 4488 4536 4494 4548
rect 6086 4536 6092 4548
rect 4488 4508 6092 4536
rect 4488 4496 4494 4508
rect 6086 4496 6092 4508
rect 6144 4496 6150 4548
rect 8110 4536 8116 4548
rect 7958 4508 8116 4536
rect 8110 4496 8116 4508
rect 8168 4496 8174 4548
rect 8861 4539 8919 4545
rect 8861 4505 8873 4539
rect 8907 4536 8919 4539
rect 9214 4536 9220 4548
rect 8907 4508 9220 4536
rect 8907 4505 8919 4508
rect 8861 4499 8919 4505
rect 9214 4496 9220 4508
rect 9272 4536 9278 4548
rect 9272 4508 16574 4536
rect 9272 4496 9278 4508
rect 16546 4480 16574 4508
rect 4246 4468 4252 4480
rect 4207 4440 4252 4468
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4338 4428 4344 4480
rect 4396 4468 4402 4480
rect 4893 4471 4951 4477
rect 4893 4468 4905 4471
rect 4396 4440 4905 4468
rect 4396 4428 4402 4440
rect 4893 4437 4905 4440
rect 4939 4437 4951 4471
rect 4893 4431 4951 4437
rect 4982 4428 4988 4480
rect 5040 4468 5046 4480
rect 6181 4471 6239 4477
rect 6181 4468 6193 4471
rect 5040 4440 6193 4468
rect 5040 4428 5046 4440
rect 6181 4437 6193 4440
rect 6227 4437 6239 4471
rect 6181 4431 6239 4437
rect 6638 4428 6644 4480
rect 6696 4468 6702 4480
rect 8662 4468 8668 4480
rect 6696 4440 8668 4468
rect 6696 4428 6702 4440
rect 8662 4428 8668 4440
rect 8720 4428 8726 4480
rect 16546 4440 16580 4480
rect 16574 4428 16580 4440
rect 16632 4428 16638 4480
rect 3036 4378 9844 4400
rect 3036 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 5194 4378
rect 5246 4326 5258 4378
rect 5310 4326 5322 4378
rect 5374 4326 9844 4378
rect 3036 4304 9844 4326
rect 3234 4224 3240 4276
rect 3292 4264 3298 4276
rect 3329 4267 3387 4273
rect 3329 4264 3341 4267
rect 3292 4236 3341 4264
rect 3292 4224 3298 4236
rect 3329 4233 3341 4236
rect 3375 4233 3387 4267
rect 5718 4264 5724 4276
rect 3329 4227 3387 4233
rect 3804 4236 5724 4264
rect 3804 4205 3832 4236
rect 5718 4224 5724 4236
rect 5776 4224 5782 4276
rect 5810 4224 5816 4276
rect 5868 4264 5874 4276
rect 5868 4236 7144 4264
rect 5868 4224 5874 4236
rect 3789 4199 3847 4205
rect 3789 4165 3801 4199
rect 3835 4165 3847 4199
rect 4062 4196 4068 4208
rect 3789 4159 3847 4165
rect 3988 4168 4068 4196
rect 3142 4088 3148 4140
rect 3200 4128 3206 4140
rect 3418 4128 3424 4140
rect 3200 4100 3424 4128
rect 3200 4088 3206 4100
rect 3418 4088 3424 4100
rect 3476 4128 3482 4140
rect 3513 4131 3571 4137
rect 3513 4128 3525 4131
rect 3476 4100 3525 4128
rect 3476 4088 3482 4100
rect 3513 4097 3525 4100
rect 3559 4097 3571 4131
rect 3513 4091 3571 4097
rect 3694 4088 3700 4140
rect 3752 4128 3758 4140
rect 3988 4137 4016 4168
rect 4062 4156 4068 4168
rect 4120 4156 4126 4208
rect 4430 4196 4436 4208
rect 4172 4168 4436 4196
rect 4172 4137 4200 4168
rect 4430 4156 4436 4168
rect 4488 4156 4494 4208
rect 5166 4156 5172 4208
rect 5224 4156 5230 4208
rect 7116 4205 7144 4236
rect 8294 4224 8300 4276
rect 8352 4264 8358 4276
rect 8757 4267 8815 4273
rect 8757 4264 8769 4267
rect 8352 4236 8769 4264
rect 8352 4224 8358 4236
rect 8757 4233 8769 4236
rect 8803 4233 8815 4267
rect 8757 4227 8815 4233
rect 9490 4224 9496 4276
rect 9548 4224 9554 4276
rect 7101 4199 7159 4205
rect 7101 4165 7113 4199
rect 7147 4165 7159 4199
rect 8018 4196 8024 4208
rect 7101 4159 7159 4165
rect 7576 4168 8024 4196
rect 3973 4131 4031 4137
rect 3973 4128 3985 4131
rect 3752 4100 3985 4128
rect 3752 4088 3758 4100
rect 3973 4097 3985 4100
rect 4019 4097 4031 4131
rect 3973 4091 4031 4097
rect 4157 4131 4215 4137
rect 4157 4097 4169 4131
rect 4203 4097 4215 4131
rect 6270 4128 6276 4140
rect 4157 4091 4215 4097
rect 4540 4100 4936 4128
rect 6231 4100 6276 4128
rect 3602 4020 3608 4072
rect 3660 4060 3666 4072
rect 4433 4063 4491 4069
rect 4433 4060 4445 4063
rect 3660 4032 4445 4060
rect 3660 4020 3666 4032
rect 4433 4029 4445 4032
rect 4479 4029 4491 4063
rect 4433 4023 4491 4029
rect 3510 3952 3516 4004
rect 3568 3992 3574 4004
rect 4540 3992 4568 4100
rect 4798 4060 4804 4072
rect 4759 4032 4804 4060
rect 4798 4020 4804 4032
rect 4856 4020 4862 4072
rect 4908 4060 4936 4100
rect 6270 4088 6276 4100
rect 6328 4088 6334 4140
rect 7190 4088 7196 4140
rect 7248 4128 7254 4140
rect 7377 4131 7435 4137
rect 7377 4128 7389 4131
rect 7248 4100 7389 4128
rect 7248 4088 7254 4100
rect 7377 4097 7389 4100
rect 7423 4097 7435 4131
rect 7377 4091 7435 4097
rect 5166 4060 5172 4072
rect 4908 4032 5172 4060
rect 5166 4020 5172 4032
rect 5224 4020 5230 4072
rect 6454 4020 6460 4072
rect 6512 4060 6518 4072
rect 7469 4063 7527 4069
rect 7469 4060 7481 4063
rect 6512 4032 7481 4060
rect 6512 4020 6518 4032
rect 7469 4029 7481 4032
rect 7515 4029 7527 4063
rect 7469 4023 7527 4029
rect 3568 3964 4568 3992
rect 3568 3952 3574 3964
rect 5902 3952 5908 4004
rect 5960 3992 5966 4004
rect 7576 3992 7604 4168
rect 8018 4156 8024 4168
rect 8076 4196 8082 4208
rect 8481 4199 8539 4205
rect 8481 4196 8493 4199
rect 8076 4168 8493 4196
rect 8076 4156 8082 4168
rect 8481 4165 8493 4168
rect 8527 4165 8539 4199
rect 8481 4159 8539 4165
rect 8570 4156 8576 4208
rect 8628 4196 8634 4208
rect 9125 4199 9183 4205
rect 9125 4196 9137 4199
rect 8628 4168 9137 4196
rect 8628 4156 8634 4168
rect 9125 4165 9137 4168
rect 9171 4196 9183 4199
rect 9508 4196 9536 4224
rect 9171 4168 9536 4196
rect 9171 4165 9183 4168
rect 9125 4159 9183 4165
rect 7653 4131 7711 4137
rect 7653 4097 7665 4131
rect 7699 4097 7711 4131
rect 7653 4091 7711 4097
rect 7668 4060 7696 4091
rect 7926 4088 7932 4140
rect 7984 4128 7990 4140
rect 8113 4131 8171 4137
rect 8113 4128 8125 4131
rect 7984 4100 8125 4128
rect 7984 4088 7990 4100
rect 8113 4097 8125 4100
rect 8159 4097 8171 4131
rect 8113 4091 8171 4097
rect 8202 4088 8208 4140
rect 8260 4128 8266 4140
rect 8662 4128 8668 4140
rect 8260 4100 8440 4128
rect 8623 4100 8668 4128
rect 8260 4088 8266 4100
rect 8297 4063 8355 4069
rect 8297 4060 8309 4063
rect 7668 4032 8309 4060
rect 8297 4029 8309 4032
rect 8343 4029 8355 4063
rect 8412 4060 8440 4100
rect 8662 4088 8668 4100
rect 8720 4088 8726 4140
rect 8938 4128 8944 4140
rect 8899 4100 8944 4128
rect 8938 4088 8944 4100
rect 8996 4088 9002 4140
rect 9493 4131 9551 4137
rect 9493 4097 9505 4131
rect 9539 4097 9551 4131
rect 9493 4091 9551 4097
rect 9508 4060 9536 4091
rect 8412 4032 9536 4060
rect 8297 4023 8355 4029
rect 5960 3964 7604 3992
rect 7837 3995 7895 4001
rect 5960 3952 5966 3964
rect 7837 3961 7849 3995
rect 7883 3992 7895 3995
rect 8202 3992 8208 4004
rect 7883 3964 8208 3992
rect 7883 3961 7895 3964
rect 7837 3955 7895 3961
rect 8202 3952 8208 3964
rect 8260 3952 8266 4004
rect 9309 3995 9367 4001
rect 9309 3992 9321 3995
rect 8312 3964 9321 3992
rect 3697 3927 3755 3933
rect 3697 3893 3709 3927
rect 3743 3924 3755 3927
rect 3878 3924 3884 3936
rect 3743 3896 3884 3924
rect 3743 3893 3755 3896
rect 3697 3887 3755 3893
rect 3878 3884 3884 3896
rect 3936 3884 3942 3936
rect 4249 3927 4307 3933
rect 4249 3893 4261 3927
rect 4295 3924 4307 3927
rect 6730 3924 6736 3936
rect 4295 3896 6736 3924
rect 4295 3893 4307 3896
rect 4249 3887 4307 3893
rect 6730 3884 6736 3896
rect 6788 3884 6794 3936
rect 6822 3884 6828 3936
rect 6880 3933 6886 3936
rect 6880 3924 6891 3933
rect 7190 3924 7196 3936
rect 6880 3896 6925 3924
rect 7151 3896 7196 3924
rect 6880 3887 6891 3896
rect 6880 3884 6886 3887
rect 7190 3884 7196 3896
rect 7248 3884 7254 3936
rect 7926 3924 7932 3936
rect 7887 3896 7932 3924
rect 7926 3884 7932 3896
rect 7984 3884 7990 3936
rect 8110 3884 8116 3936
rect 8168 3924 8174 3936
rect 8312 3924 8340 3964
rect 9309 3961 9321 3964
rect 9355 3961 9367 3995
rect 9309 3955 9367 3961
rect 8168 3896 8340 3924
rect 8168 3884 8174 3896
rect 3036 3834 9844 3856
rect 3036 3782 7566 3834
rect 7618 3782 7630 3834
rect 7682 3782 7694 3834
rect 7746 3782 7758 3834
rect 7810 3782 7822 3834
rect 7874 3782 9844 3834
rect 3036 3760 9844 3782
rect 3602 3720 3608 3732
rect 3563 3692 3608 3720
rect 3602 3680 3608 3692
rect 3660 3680 3666 3732
rect 5166 3680 5172 3732
rect 5224 3720 5230 3732
rect 5353 3723 5411 3729
rect 5353 3720 5365 3723
rect 5224 3692 5365 3720
rect 5224 3680 5230 3692
rect 5353 3689 5365 3692
rect 5399 3689 5411 3723
rect 5353 3683 5411 3689
rect 6273 3723 6331 3729
rect 6273 3689 6285 3723
rect 6319 3720 6331 3723
rect 6362 3720 6368 3732
rect 6319 3692 6368 3720
rect 6319 3689 6331 3692
rect 6273 3683 6331 3689
rect 6362 3680 6368 3692
rect 6420 3720 6426 3732
rect 6638 3720 6644 3732
rect 6420 3692 6644 3720
rect 6420 3680 6426 3692
rect 6638 3680 6644 3692
rect 6696 3680 6702 3732
rect 6730 3680 6736 3732
rect 6788 3720 6794 3732
rect 6788 3692 8340 3720
rect 6788 3680 6794 3692
rect 3418 3612 3424 3664
rect 3476 3652 3482 3664
rect 4614 3652 4620 3664
rect 3476 3624 4620 3652
rect 3476 3612 3482 3624
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 4709 3655 4767 3661
rect 4709 3621 4721 3655
rect 4755 3652 4767 3655
rect 5534 3652 5540 3664
rect 4755 3624 5540 3652
rect 4755 3621 4767 3624
rect 4709 3615 4767 3621
rect 5534 3612 5540 3624
rect 5592 3612 5598 3664
rect 5166 3584 5172 3596
rect 4540 3556 5172 3584
rect 3418 3516 3424 3528
rect 3379 3488 3424 3516
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3697 3519 3755 3525
rect 3697 3485 3709 3519
rect 3743 3516 3755 3519
rect 3973 3519 4031 3525
rect 3973 3516 3985 3519
rect 3743 3488 3985 3516
rect 3743 3485 3755 3488
rect 3697 3479 3755 3485
rect 3973 3485 3985 3488
rect 4019 3516 4031 3519
rect 4154 3516 4160 3528
rect 4019 3488 4160 3516
rect 4019 3485 4031 3488
rect 3973 3479 4031 3485
rect 4154 3476 4160 3488
rect 4212 3476 4218 3528
rect 4246 3476 4252 3528
rect 4304 3516 4310 3528
rect 4540 3525 4568 3556
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 7190 3584 7196 3596
rect 5276 3556 7196 3584
rect 4525 3519 4583 3525
rect 4304 3488 4349 3516
rect 4304 3476 4310 3488
rect 4525 3485 4537 3519
rect 4571 3485 4583 3519
rect 4525 3479 4583 3485
rect 4890 3476 4896 3528
rect 4948 3476 4954 3528
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5276 3516 5304 3556
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 5031 3488 5304 3516
rect 5721 3519 5779 3525
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 5721 3485 5733 3519
rect 5767 3516 5779 3519
rect 5994 3516 6000 3528
rect 5767 3488 6000 3516
rect 5767 3485 5779 3488
rect 5721 3479 5779 3485
rect 5994 3476 6000 3488
rect 6052 3476 6058 3528
rect 6365 3519 6423 3525
rect 6365 3485 6377 3519
rect 6411 3485 6423 3519
rect 6730 3516 6736 3528
rect 6691 3488 6736 3516
rect 6365 3479 6423 3485
rect 4908 3448 4936 3476
rect 5074 3448 5080 3460
rect 4908 3420 5080 3448
rect 5074 3408 5080 3420
rect 5132 3408 5138 3460
rect 5261 3451 5319 3457
rect 5261 3417 5273 3451
rect 5307 3448 5319 3451
rect 5902 3448 5908 3460
rect 5307 3420 5908 3448
rect 5307 3417 5319 3420
rect 5261 3411 5319 3417
rect 5902 3408 5908 3420
rect 5960 3408 5966 3460
rect 6086 3448 6092 3460
rect 6047 3420 6092 3448
rect 6086 3408 6092 3420
rect 6144 3408 6150 3460
rect 3694 3340 3700 3392
rect 3752 3380 3758 3392
rect 3881 3383 3939 3389
rect 3881 3380 3893 3383
rect 3752 3352 3893 3380
rect 3752 3340 3758 3352
rect 3881 3349 3893 3352
rect 3927 3349 3939 3383
rect 3881 3343 3939 3349
rect 4157 3383 4215 3389
rect 4157 3349 4169 3383
rect 4203 3380 4215 3383
rect 4246 3380 4252 3392
rect 4203 3352 4252 3380
rect 4203 3349 4215 3352
rect 4157 3343 4215 3349
rect 4246 3340 4252 3352
rect 4304 3340 4310 3392
rect 4430 3380 4436 3392
rect 4391 3352 4436 3380
rect 4430 3340 4436 3352
rect 4488 3340 4494 3392
rect 4893 3383 4951 3389
rect 4893 3349 4905 3383
rect 4939 3380 4951 3383
rect 6380 3380 6408 3479
rect 6730 3476 6736 3488
rect 6788 3476 6794 3528
rect 8202 3516 8208 3528
rect 8163 3488 8208 3516
rect 8202 3476 8208 3488
rect 8260 3476 8266 3528
rect 8312 3516 8340 3692
rect 8754 3680 8760 3732
rect 8812 3729 8818 3732
rect 8812 3720 8823 3729
rect 9493 3723 9551 3729
rect 8812 3692 8857 3720
rect 8812 3683 8823 3692
rect 9493 3689 9505 3723
rect 9539 3720 9551 3723
rect 9582 3720 9588 3732
rect 9539 3692 9588 3720
rect 9539 3689 9551 3692
rect 9493 3683 9551 3689
rect 8812 3680 8818 3683
rect 9582 3680 9588 3692
rect 9640 3680 9646 3732
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8312 3488 9137 3516
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 7926 3448 7932 3460
rect 7866 3420 7932 3448
rect 7926 3408 7932 3420
rect 7984 3408 7990 3460
rect 9217 3451 9275 3457
rect 9217 3448 9229 3451
rect 8036 3420 9229 3448
rect 4939 3352 6408 3380
rect 4939 3349 4951 3352
rect 4893 3343 4951 3349
rect 6730 3340 6736 3392
rect 6788 3380 6794 3392
rect 7006 3380 7012 3392
rect 6788 3352 7012 3380
rect 6788 3340 6794 3352
rect 7006 3340 7012 3352
rect 7064 3340 7070 3392
rect 7374 3340 7380 3392
rect 7432 3380 7438 3392
rect 8036 3380 8064 3420
rect 9217 3417 9229 3420
rect 9263 3417 9275 3451
rect 9217 3411 9275 3417
rect 8938 3380 8944 3392
rect 7432 3352 8064 3380
rect 8899 3352 8944 3380
rect 7432 3340 7438 3352
rect 8938 3340 8944 3352
rect 8996 3340 9002 3392
rect 3036 3290 9844 3312
rect 3036 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 5194 3290
rect 5246 3238 5258 3290
rect 5310 3238 5322 3290
rect 5374 3238 9844 3290
rect 3036 3216 9844 3238
rect 3602 3136 3608 3188
rect 3660 3176 3666 3188
rect 3878 3176 3884 3188
rect 3660 3148 3884 3176
rect 3660 3136 3666 3148
rect 3878 3136 3884 3148
rect 3936 3176 3942 3188
rect 3936 3148 6316 3176
rect 3936 3136 3942 3148
rect 4430 3068 4436 3120
rect 4488 3068 4494 3120
rect 3421 3043 3479 3049
rect 3421 3009 3433 3043
rect 3467 3009 3479 3043
rect 3694 3040 3700 3052
rect 3655 3012 3700 3040
rect 3421 3003 3479 3009
rect 3436 2972 3464 3003
rect 3694 3000 3700 3012
rect 3752 3000 3758 3052
rect 5534 3040 5540 3052
rect 3804 3012 4200 3040
rect 5495 3012 5540 3040
rect 3804 2972 3832 3012
rect 4062 2972 4068 2984
rect 3436 2944 3832 2972
rect 4023 2944 4068 2972
rect 4062 2932 4068 2944
rect 4120 2932 4126 2984
rect 4172 2972 4200 3012
rect 5534 3000 5540 3012
rect 5592 3000 5598 3052
rect 6288 3049 6316 3148
rect 6362 3136 6368 3188
rect 6420 3176 6426 3188
rect 7374 3176 7380 3188
rect 6420 3148 7380 3176
rect 6420 3136 6426 3148
rect 7374 3136 7380 3148
rect 7432 3136 7438 3188
rect 8021 3179 8079 3185
rect 8021 3145 8033 3179
rect 8067 3145 8079 3179
rect 8021 3139 8079 3145
rect 8297 3179 8355 3185
rect 8297 3145 8309 3179
rect 8343 3176 8355 3179
rect 8478 3176 8484 3188
rect 8343 3148 8484 3176
rect 8343 3145 8355 3148
rect 8297 3139 8355 3145
rect 6454 3068 6460 3120
rect 6512 3108 6518 3120
rect 6549 3111 6607 3117
rect 6549 3108 6561 3111
rect 6512 3080 6561 3108
rect 6512 3068 6518 3080
rect 6549 3077 6561 3080
rect 6595 3077 6607 3111
rect 6549 3071 6607 3077
rect 7006 3068 7012 3120
rect 7064 3068 7070 3120
rect 8036 3108 8064 3139
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 8386 3108 8392 3120
rect 8036 3080 8392 3108
rect 8386 3068 8392 3080
rect 8444 3108 8450 3120
rect 8444 3080 8984 3108
rect 8444 3068 8450 3080
rect 8956 3049 8984 3080
rect 6273 3043 6331 3049
rect 6273 3009 6285 3043
rect 6319 3009 6331 3043
rect 6273 3003 6331 3009
rect 8941 3043 8999 3049
rect 8941 3009 8953 3043
rect 8987 3009 8999 3043
rect 8941 3003 8999 3009
rect 9033 3043 9091 3049
rect 9033 3009 9045 3043
rect 9079 3040 9091 3043
rect 9306 3040 9312 3052
rect 9079 3012 9312 3040
rect 9079 3009 9091 3012
rect 9033 3003 9091 3009
rect 9306 3000 9312 3012
rect 9364 3000 9370 3052
rect 9493 3043 9551 3049
rect 9493 3009 9505 3043
rect 9539 3040 9551 3043
rect 9582 3040 9588 3052
rect 9539 3012 9588 3040
rect 9539 3009 9551 3012
rect 9493 3003 9551 3009
rect 9582 3000 9588 3012
rect 9640 3000 9646 3052
rect 4338 2972 4344 2984
rect 4172 2944 4344 2972
rect 4338 2932 4344 2944
rect 4396 2932 4402 2984
rect 6638 2972 6644 2984
rect 6012 2944 6644 2972
rect 3510 2864 3516 2916
rect 3568 2904 3574 2916
rect 3605 2907 3663 2913
rect 3605 2904 3617 2907
rect 3568 2876 3617 2904
rect 3568 2864 3574 2876
rect 3605 2873 3617 2876
rect 3651 2873 3663 2907
rect 3605 2867 3663 2873
rect 4062 2796 4068 2848
rect 4120 2836 4126 2848
rect 6012 2836 6040 2944
rect 6638 2932 6644 2944
rect 6696 2932 6702 2984
rect 8478 2864 8484 2916
rect 8536 2904 8542 2916
rect 9401 2907 9459 2913
rect 9401 2904 9413 2907
rect 8536 2876 9413 2904
rect 8536 2864 8542 2876
rect 9401 2873 9413 2876
rect 9447 2873 9459 2907
rect 9401 2867 9459 2873
rect 4120 2808 6040 2836
rect 6101 2839 6159 2845
rect 4120 2796 4126 2808
rect 6101 2805 6113 2839
rect 6147 2836 6159 2839
rect 6546 2836 6552 2848
rect 6147 2808 6552 2836
rect 6147 2805 6159 2808
rect 6101 2799 6159 2805
rect 6546 2796 6552 2808
rect 6604 2796 6610 2848
rect 9214 2836 9220 2848
rect 9175 2808 9220 2836
rect 9214 2796 9220 2808
rect 9272 2796 9278 2848
rect 3036 2746 9844 2768
rect 3036 2694 7566 2746
rect 7618 2694 7630 2746
rect 7682 2694 7694 2746
rect 7746 2694 7758 2746
rect 7810 2694 7822 2746
rect 7874 2694 9844 2746
rect 3036 2672 9844 2694
rect 4246 2592 4252 2644
rect 4304 2632 4310 2644
rect 4614 2632 4620 2644
rect 4304 2604 4620 2632
rect 4304 2592 4310 2604
rect 4614 2592 4620 2604
rect 4672 2632 4678 2644
rect 5442 2632 5448 2644
rect 4672 2604 5448 2632
rect 4672 2592 4678 2604
rect 5442 2592 5448 2604
rect 5500 2592 5506 2644
rect 5905 2635 5963 2641
rect 5905 2601 5917 2635
rect 5951 2632 5963 2635
rect 6270 2632 6276 2644
rect 5951 2604 6276 2632
rect 5951 2601 5963 2604
rect 5905 2595 5963 2601
rect 6270 2592 6276 2604
rect 6328 2592 6334 2644
rect 8386 2592 8392 2644
rect 8444 2641 8450 2644
rect 8444 2632 8455 2641
rect 8444 2604 8489 2632
rect 8444 2595 8455 2604
rect 8444 2592 8450 2595
rect 5460 2564 5488 2592
rect 5460 2536 6144 2564
rect 3602 2496 3608 2508
rect 3344 2468 3608 2496
rect 3344 2440 3372 2468
rect 3602 2456 3608 2468
rect 3660 2456 3666 2508
rect 4154 2456 4160 2508
rect 4212 2496 4218 2508
rect 5445 2499 5503 2505
rect 4212 2468 5396 2496
rect 4212 2456 4218 2468
rect 3326 2428 3332 2440
rect 3287 2400 3332 2428
rect 3326 2388 3332 2400
rect 3384 2388 3390 2440
rect 5368 2437 5396 2468
rect 5445 2465 5457 2499
rect 5491 2496 5503 2499
rect 5997 2499 6055 2505
rect 5997 2496 6009 2499
rect 5491 2468 6009 2496
rect 5491 2465 5503 2468
rect 5445 2459 5503 2465
rect 5997 2465 6009 2468
rect 6043 2465 6055 2499
rect 6116 2496 6144 2536
rect 7006 2496 7012 2508
rect 6116 2468 7012 2496
rect 5997 2459 6055 2465
rect 7006 2456 7012 2468
rect 7064 2456 7070 2508
rect 8938 2496 8944 2508
rect 7852 2468 8944 2496
rect 5353 2431 5411 2437
rect 5353 2397 5365 2431
rect 5399 2397 5411 2431
rect 5353 2391 5411 2397
rect 5721 2431 5779 2437
rect 5721 2397 5733 2431
rect 5767 2428 5779 2431
rect 5902 2428 5908 2440
rect 5767 2400 5908 2428
rect 5767 2397 5779 2400
rect 5721 2391 5779 2397
rect 5902 2388 5908 2400
rect 5960 2388 5966 2440
rect 6362 2428 6368 2440
rect 6323 2400 6368 2428
rect 6362 2388 6368 2400
rect 6420 2388 6426 2440
rect 7852 2437 7880 2468
rect 8938 2456 8944 2468
rect 8996 2456 9002 2508
rect 9033 2499 9091 2505
rect 9033 2465 9045 2499
rect 9079 2496 9091 2499
rect 9122 2496 9128 2508
rect 9079 2468 9128 2496
rect 9079 2465 9091 2468
rect 9033 2459 9091 2465
rect 9122 2456 9128 2468
rect 9180 2456 9186 2508
rect 7837 2431 7895 2437
rect 7837 2397 7849 2431
rect 7883 2397 7895 2431
rect 7837 2391 7895 2397
rect 3605 2363 3663 2369
rect 3605 2329 3617 2363
rect 3651 2329 3663 2363
rect 3605 2323 3663 2329
rect 3620 2292 3648 2323
rect 4246 2320 4252 2372
rect 4304 2320 4310 2372
rect 6730 2320 6736 2372
rect 6788 2320 6794 2372
rect 9214 2360 9220 2372
rect 9175 2332 9220 2360
rect 9214 2320 9220 2332
rect 9272 2320 9278 2372
rect 9306 2320 9312 2372
rect 9364 2360 9370 2372
rect 9582 2360 9588 2372
rect 9364 2332 9588 2360
rect 9364 2320 9370 2332
rect 9582 2320 9588 2332
rect 9640 2320 9646 2372
rect 4614 2292 4620 2304
rect 3620 2264 4620 2292
rect 4614 2252 4620 2264
rect 4672 2252 4678 2304
rect 5077 2295 5135 2301
rect 5077 2261 5089 2295
rect 5123 2292 5135 2295
rect 5442 2292 5448 2304
rect 5123 2264 5448 2292
rect 5123 2261 5135 2264
rect 5077 2255 5135 2261
rect 5442 2252 5448 2264
rect 5500 2252 5506 2304
rect 3036 2202 9844 2224
rect 3036 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 5194 2202
rect 5246 2150 5258 2202
rect 5310 2150 5322 2202
rect 5374 2150 9844 2202
rect 3036 2128 9844 2150
rect 2682 2048 2688 2100
rect 2740 2088 2746 2100
rect 2740 2060 6592 2088
rect 2740 2048 2746 2060
rect 3513 2023 3571 2029
rect 3513 1989 3525 2023
rect 3559 2020 3571 2023
rect 3697 2023 3755 2029
rect 3697 2020 3709 2023
rect 3559 1992 3709 2020
rect 3559 1989 3571 1992
rect 3513 1983 3571 1989
rect 3697 1989 3709 1992
rect 3743 2020 3755 2023
rect 3786 2020 3792 2032
rect 3743 1992 3792 2020
rect 3743 1989 3755 1992
rect 3697 1983 3755 1989
rect 3786 1980 3792 1992
rect 3844 1980 3850 2032
rect 3881 2023 3939 2029
rect 3881 1989 3893 2023
rect 3927 2020 3939 2023
rect 4341 2023 4399 2029
rect 4341 2020 4353 2023
rect 3927 1992 4353 2020
rect 3927 1989 3939 1992
rect 3881 1983 3939 1989
rect 4341 1989 4353 1992
rect 4387 2020 4399 2023
rect 4522 2020 4528 2032
rect 4387 1992 4528 2020
rect 4387 1989 4399 1992
rect 4341 1983 4399 1989
rect 4522 1980 4528 1992
rect 4580 1980 4586 2032
rect 5534 1980 5540 2032
rect 5592 1980 5598 2032
rect 3326 1912 3332 1964
rect 3384 1952 3390 1964
rect 6564 1961 6592 2060
rect 7282 2048 7288 2100
rect 7340 2088 7346 2100
rect 8297 2091 8355 2097
rect 8297 2088 8309 2091
rect 7340 2060 8309 2088
rect 7340 2048 7346 2060
rect 8297 2057 8309 2060
rect 8343 2057 8355 2091
rect 8297 2051 8355 2057
rect 8573 2091 8631 2097
rect 8573 2057 8585 2091
rect 8619 2088 8631 2091
rect 8662 2088 8668 2100
rect 8619 2060 8668 2088
rect 8619 2057 8631 2060
rect 8573 2051 8631 2057
rect 8662 2048 8668 2060
rect 8720 2048 8726 2100
rect 9030 2088 9036 2100
rect 8991 2060 9036 2088
rect 9030 2048 9036 2060
rect 9088 2048 9094 2100
rect 4617 1955 4675 1961
rect 4617 1952 4629 1955
rect 3384 1924 4629 1952
rect 3384 1912 3390 1924
rect 4617 1921 4629 1924
rect 4663 1921 4675 1955
rect 4617 1915 4675 1921
rect 6549 1955 6607 1961
rect 6549 1921 6561 1955
rect 6595 1921 6607 1955
rect 6549 1915 6607 1921
rect 8113 1955 8171 1961
rect 8113 1921 8125 1955
rect 8159 1952 8171 1955
rect 8478 1952 8484 1964
rect 8159 1924 8484 1952
rect 8159 1921 8171 1924
rect 8113 1915 8171 1921
rect 8478 1912 8484 1924
rect 8536 1912 8542 1964
rect 8849 1955 8907 1961
rect 8849 1921 8861 1955
rect 8895 1952 8907 1955
rect 8941 1955 8999 1961
rect 8941 1952 8953 1955
rect 8895 1924 8953 1952
rect 8895 1921 8907 1924
rect 8849 1915 8907 1921
rect 8941 1921 8953 1924
rect 8987 1952 8999 1955
rect 16574 1952 16580 1964
rect 8987 1924 16580 1952
rect 8987 1921 8999 1924
rect 8941 1915 8999 1921
rect 16574 1912 16580 1924
rect 16632 1912 16638 1964
rect 4893 1887 4951 1893
rect 4893 1853 4905 1887
rect 4939 1884 4951 1887
rect 5442 1884 5448 1896
rect 4939 1856 5448 1884
rect 4939 1853 4951 1856
rect 4893 1847 4951 1853
rect 5442 1844 5448 1856
rect 5500 1844 5506 1896
rect 6365 1887 6423 1893
rect 6365 1853 6377 1887
rect 6411 1884 6423 1887
rect 6454 1884 6460 1896
rect 6411 1856 6460 1884
rect 6411 1853 6423 1856
rect 6365 1847 6423 1853
rect 6454 1844 6460 1856
rect 6512 1844 6518 1896
rect 9398 1884 9404 1896
rect 9359 1856 9404 1884
rect 9398 1844 9404 1856
rect 9456 1844 9462 1896
rect 8021 1819 8079 1825
rect 8021 1785 8033 1819
rect 8067 1816 8079 1819
rect 20622 1816 20628 1828
rect 8067 1788 20628 1816
rect 8067 1785 8079 1788
rect 8021 1779 8079 1785
rect 20622 1776 20628 1788
rect 20680 1776 20686 1828
rect 4065 1751 4123 1757
rect 4065 1717 4077 1751
rect 4111 1748 4123 1751
rect 4433 1751 4491 1757
rect 4433 1748 4445 1751
rect 4111 1720 4445 1748
rect 4111 1717 4123 1720
rect 4065 1711 4123 1717
rect 4433 1717 4445 1720
rect 4479 1748 4491 1751
rect 4890 1748 4896 1760
rect 4479 1720 4896 1748
rect 4479 1717 4491 1720
rect 4433 1711 4491 1717
rect 4890 1708 4896 1720
rect 4948 1708 4954 1760
rect 9214 1748 9220 1760
rect 9175 1720 9220 1748
rect 9214 1708 9220 1720
rect 9272 1708 9278 1760
rect 3036 1658 9844 1680
rect 3036 1606 7566 1658
rect 7618 1606 7630 1658
rect 7682 1606 7694 1658
rect 7746 1606 7758 1658
rect 7810 1606 7822 1658
rect 7874 1606 9844 1658
rect 3036 1584 9844 1606
rect 4614 1504 4620 1556
rect 4672 1544 4678 1556
rect 5077 1547 5135 1553
rect 5077 1544 5089 1547
rect 4672 1516 5089 1544
rect 4672 1504 4678 1516
rect 5077 1513 5089 1516
rect 5123 1513 5135 1547
rect 5077 1507 5135 1513
rect 3326 1408 3332 1420
rect 3287 1380 3332 1408
rect 3326 1368 3332 1380
rect 3384 1368 3390 1420
rect 3605 1411 3663 1417
rect 3605 1377 3617 1411
rect 3651 1408 3663 1411
rect 3970 1408 3976 1420
rect 3651 1380 3976 1408
rect 3651 1377 3663 1380
rect 3605 1371 3663 1377
rect 3970 1368 3976 1380
rect 4028 1368 4034 1420
rect 5092 1408 5120 1507
rect 6362 1504 6368 1556
rect 6420 1544 6426 1556
rect 6457 1547 6515 1553
rect 6457 1544 6469 1547
rect 6420 1516 6469 1544
rect 6420 1504 6426 1516
rect 6457 1513 6469 1516
rect 6503 1513 6515 1547
rect 6457 1507 6515 1513
rect 8021 1547 8079 1553
rect 8021 1513 8033 1547
rect 8067 1544 8079 1547
rect 8662 1544 8668 1556
rect 8067 1516 8668 1544
rect 8067 1513 8079 1516
rect 8021 1507 8079 1513
rect 8662 1504 8668 1516
rect 8720 1504 8726 1556
rect 9217 1547 9275 1553
rect 9217 1513 9229 1547
rect 9263 1544 9275 1547
rect 9306 1544 9312 1556
rect 9263 1516 9312 1544
rect 9263 1513 9275 1516
rect 9217 1507 9275 1513
rect 9306 1504 9312 1516
rect 9364 1504 9370 1556
rect 5537 1479 5595 1485
rect 5537 1445 5549 1479
rect 5583 1476 5595 1479
rect 6730 1476 6736 1488
rect 5583 1448 6736 1476
rect 5583 1445 5595 1448
rect 5537 1439 5595 1445
rect 6730 1436 6736 1448
rect 6788 1436 6794 1488
rect 5092 1380 5856 1408
rect 4982 1300 4988 1352
rect 5040 1340 5046 1352
rect 5353 1343 5411 1349
rect 5353 1340 5365 1343
rect 5040 1312 5365 1340
rect 5040 1300 5046 1312
rect 5353 1309 5365 1312
rect 5399 1309 5411 1343
rect 5353 1303 5411 1309
rect 5442 1300 5448 1352
rect 5500 1340 5506 1352
rect 5721 1343 5779 1349
rect 5721 1340 5733 1343
rect 5500 1312 5733 1340
rect 5500 1300 5506 1312
rect 5721 1309 5733 1312
rect 5767 1309 5779 1343
rect 5828 1340 5856 1380
rect 6380 1380 7236 1408
rect 6380 1340 6408 1380
rect 5828 1312 6408 1340
rect 5721 1303 5779 1309
rect 6454 1300 6460 1352
rect 6512 1340 6518 1352
rect 7208 1349 7236 1380
rect 7101 1343 7159 1349
rect 7101 1340 7113 1343
rect 6512 1312 7113 1340
rect 6512 1300 6518 1312
rect 7101 1309 7113 1312
rect 7147 1309 7159 1343
rect 7101 1303 7159 1309
rect 7193 1343 7251 1349
rect 7193 1309 7205 1343
rect 7239 1309 7251 1343
rect 7193 1303 7251 1309
rect 4246 1232 4252 1284
rect 4304 1232 4310 1284
rect 4890 1232 4896 1284
rect 4948 1272 4954 1284
rect 6365 1275 6423 1281
rect 6365 1272 6377 1275
rect 4948 1244 6377 1272
rect 4948 1232 4954 1244
rect 6365 1241 6377 1244
rect 6411 1241 6423 1275
rect 6365 1235 6423 1241
rect 6638 1232 6644 1284
rect 6696 1272 6702 1284
rect 7837 1275 7895 1281
rect 7837 1272 7849 1275
rect 6696 1244 7849 1272
rect 6696 1232 6702 1244
rect 7837 1241 7849 1244
rect 7883 1241 7895 1275
rect 7837 1235 7895 1241
rect 7006 1164 7012 1216
rect 7064 1204 7070 1216
rect 8297 1207 8355 1213
rect 8297 1204 8309 1207
rect 7064 1176 8309 1204
rect 7064 1164 7070 1176
rect 8297 1173 8309 1176
rect 8343 1204 8355 1207
rect 8481 1207 8539 1213
rect 8481 1204 8493 1207
rect 8343 1176 8493 1204
rect 8343 1173 8355 1176
rect 8297 1167 8355 1173
rect 8481 1173 8493 1176
rect 8527 1204 8539 1207
rect 8665 1207 8723 1213
rect 8665 1204 8677 1207
rect 8527 1176 8677 1204
rect 8527 1173 8539 1176
rect 8481 1167 8539 1173
rect 8665 1173 8677 1176
rect 8711 1204 8723 1207
rect 8849 1207 8907 1213
rect 8849 1204 8861 1207
rect 8711 1176 8861 1204
rect 8711 1173 8723 1176
rect 8665 1167 8723 1173
rect 8849 1173 8861 1176
rect 8895 1204 8907 1207
rect 9309 1207 9367 1213
rect 9309 1204 9321 1207
rect 8895 1176 9321 1204
rect 8895 1173 8907 1176
rect 8849 1167 8907 1173
rect 9309 1173 9321 1176
rect 9355 1173 9367 1207
rect 9309 1167 9367 1173
rect 3036 1114 9844 1136
rect 3036 1062 5066 1114
rect 5118 1062 5130 1114
rect 5182 1062 5194 1114
rect 5246 1062 5258 1114
rect 5310 1062 5322 1114
rect 5374 1062 9844 1114
rect 3036 1040 9844 1062
<< via1 >>
rect 2780 11568 2832 11620
rect 4252 11568 4304 11620
rect 1860 11500 1912 11552
rect 4988 11500 5040 11552
rect 2566 11398 2618 11450
rect 2630 11398 2682 11450
rect 2694 11398 2746 11450
rect 2758 11398 2810 11450
rect 2822 11398 2874 11450
rect 7566 11398 7618 11450
rect 7630 11398 7682 11450
rect 7694 11398 7746 11450
rect 7758 11398 7810 11450
rect 7822 11398 7874 11450
rect 1400 11296 1452 11348
rect 2412 11296 2464 11348
rect 1860 11228 1912 11280
rect 2320 11228 2372 11280
rect 2964 11228 3016 11280
rect 3516 11228 3568 11280
rect 4620 11296 4672 11348
rect 5448 11296 5500 11348
rect 5632 11296 5684 11348
rect 8116 11296 8168 11348
rect 8668 11296 8720 11348
rect 4528 11271 4580 11280
rect 4528 11237 4537 11271
rect 4537 11237 4571 11271
rect 4571 11237 4580 11271
rect 4528 11228 4580 11237
rect 5080 11228 5132 11280
rect 4620 11203 4672 11212
rect 1676 11092 1728 11144
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 2688 11092 2740 11144
rect 4620 11169 4629 11203
rect 4629 11169 4663 11203
rect 4663 11169 4672 11203
rect 4620 11160 4672 11169
rect 5908 11160 5960 11212
rect 7932 11228 7984 11280
rect 16580 11228 16632 11280
rect 7104 11160 7156 11212
rect 4344 11135 4396 11144
rect 4344 11101 4353 11135
rect 4353 11101 4387 11135
rect 4387 11101 4396 11135
rect 4344 11092 4396 11101
rect 6092 11092 6144 11144
rect 6184 11135 6236 11144
rect 6184 11101 6193 11135
rect 6193 11101 6227 11135
rect 6227 11101 6236 11135
rect 6184 11092 6236 11101
rect 6460 11092 6512 11144
rect 7196 11135 7248 11144
rect 7196 11101 7205 11135
rect 7205 11101 7239 11135
rect 7239 11101 7248 11135
rect 7196 11092 7248 11101
rect 7564 11092 7616 11144
rect 1952 10999 2004 11008
rect 1952 10965 1961 10999
rect 1961 10965 1995 10999
rect 1995 10965 2004 10999
rect 1952 10956 2004 10965
rect 2136 10956 2188 11008
rect 2964 11024 3016 11076
rect 3056 11067 3108 11076
rect 3056 11033 3065 11067
rect 3065 11033 3099 11067
rect 3099 11033 3108 11067
rect 3240 11067 3292 11076
rect 3056 11024 3108 11033
rect 3240 11033 3249 11067
rect 3249 11033 3283 11067
rect 3283 11033 3292 11067
rect 3240 11024 3292 11033
rect 3424 11024 3476 11076
rect 5448 11067 5500 11076
rect 5448 11033 5457 11067
rect 5457 11033 5491 11067
rect 5491 11033 5500 11067
rect 5448 11024 5500 11033
rect 5724 11024 5776 11076
rect 6920 11067 6972 11076
rect 6920 11033 6929 11067
rect 6929 11033 6963 11067
rect 6963 11033 6972 11067
rect 6920 11024 6972 11033
rect 7012 11024 7064 11076
rect 7380 11024 7432 11076
rect 8024 11067 8076 11076
rect 8024 11033 8033 11067
rect 8033 11033 8067 11067
rect 8067 11033 8076 11067
rect 8024 11024 8076 11033
rect 3608 10956 3660 11008
rect 4896 10999 4948 11008
rect 4896 10965 4905 10999
rect 4905 10965 4939 10999
rect 4939 10965 4948 10999
rect 4896 10956 4948 10965
rect 6184 10956 6236 11008
rect 7840 10956 7892 11008
rect 8392 10999 8444 11008
rect 8392 10965 8401 10999
rect 8401 10965 8435 10999
rect 8435 10965 8444 10999
rect 8392 10956 8444 10965
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 5194 10854 5246 10906
rect 5258 10854 5310 10906
rect 5322 10854 5374 10906
rect 4344 10752 4396 10804
rect 1676 10727 1728 10736
rect 1676 10693 1685 10727
rect 1685 10693 1719 10727
rect 1719 10693 1728 10727
rect 1676 10684 1728 10693
rect 3240 10684 3292 10736
rect 1492 10659 1544 10668
rect 1492 10625 1501 10659
rect 1501 10625 1535 10659
rect 1535 10625 1544 10659
rect 1492 10616 1544 10625
rect 1952 10616 2004 10668
rect 3608 10659 3660 10668
rect 3608 10625 3617 10659
rect 3617 10625 3651 10659
rect 3651 10625 3660 10659
rect 3608 10616 3660 10625
rect 4620 10616 4672 10668
rect 5448 10752 5500 10804
rect 7840 10795 7892 10804
rect 6092 10684 6144 10736
rect 7840 10761 7849 10795
rect 7849 10761 7883 10795
rect 7883 10761 7892 10795
rect 7840 10752 7892 10761
rect 5540 10616 5592 10668
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 1860 10548 1912 10600
rect 2136 10591 2188 10600
rect 2136 10557 2145 10591
rect 2145 10557 2179 10591
rect 2179 10557 2188 10591
rect 2136 10548 2188 10557
rect 6736 10616 6788 10668
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 8116 10616 8168 10668
rect 9312 10659 9364 10668
rect 9312 10625 9321 10659
rect 9321 10625 9355 10659
rect 9355 10625 9364 10659
rect 9312 10616 9364 10625
rect 4804 10455 4856 10464
rect 4804 10421 4813 10455
rect 4813 10421 4847 10455
rect 4847 10421 4856 10455
rect 4804 10412 4856 10421
rect 5816 10455 5868 10464
rect 5816 10421 5825 10455
rect 5825 10421 5859 10455
rect 5859 10421 5868 10455
rect 5816 10412 5868 10421
rect 8392 10548 8444 10600
rect 7564 10480 7616 10532
rect 7104 10412 7156 10464
rect 7288 10455 7340 10464
rect 7288 10421 7297 10455
rect 7297 10421 7331 10455
rect 7331 10421 7340 10455
rect 7288 10412 7340 10421
rect 7472 10455 7524 10464
rect 7472 10421 7481 10455
rect 7481 10421 7515 10455
rect 7515 10421 7524 10455
rect 7472 10412 7524 10421
rect 8116 10455 8168 10464
rect 8116 10421 8125 10455
rect 8125 10421 8159 10455
rect 8159 10421 8168 10455
rect 8116 10412 8168 10421
rect 8300 10412 8352 10464
rect 16580 10412 16632 10464
rect 2566 10310 2618 10362
rect 2630 10310 2682 10362
rect 2694 10310 2746 10362
rect 2758 10310 2810 10362
rect 2822 10310 2874 10362
rect 7566 10310 7618 10362
rect 7630 10310 7682 10362
rect 7694 10310 7746 10362
rect 7758 10310 7810 10362
rect 7822 10310 7874 10362
rect 1492 10208 1544 10260
rect 6736 10208 6788 10260
rect 7196 10208 7248 10260
rect 2136 10140 2188 10192
rect 3240 10140 3292 10192
rect 8208 10140 8260 10192
rect 7288 10072 7340 10124
rect 3056 10004 3108 10056
rect 3792 10047 3844 10056
rect 3792 10013 3801 10047
rect 3801 10013 3835 10047
rect 3835 10013 3844 10047
rect 3792 10004 3844 10013
rect 4896 10004 4948 10056
rect 6184 10004 6236 10056
rect 8484 10004 8536 10056
rect 9496 10072 9548 10124
rect 9404 10047 9456 10056
rect 9404 10013 9413 10047
rect 9413 10013 9447 10047
rect 9447 10013 9456 10047
rect 9404 10004 9456 10013
rect 7472 9936 7524 9988
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 5194 9766 5246 9818
rect 5258 9766 5310 9818
rect 5322 9766 5374 9818
rect 1860 9664 1912 9716
rect 7288 9664 7340 9716
rect 8208 9664 8260 9716
rect 9496 9707 9548 9716
rect 9496 9673 9505 9707
rect 9505 9673 9539 9707
rect 9539 9673 9548 9707
rect 9496 9664 9548 9673
rect 16672 9664 16724 9716
rect 1492 9639 1544 9648
rect 1492 9605 1501 9639
rect 1501 9605 1535 9639
rect 1535 9605 1544 9639
rect 1492 9596 1544 9605
rect 4528 9596 4580 9648
rect 7932 9596 7984 9648
rect 3148 9528 3200 9580
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 5816 9528 5868 9580
rect 6276 9528 6328 9580
rect 6552 9571 6604 9580
rect 6552 9537 6561 9571
rect 6561 9537 6595 9571
rect 6595 9537 6604 9571
rect 6552 9528 6604 9537
rect 7012 9528 7064 9580
rect 8116 9528 8168 9580
rect 4068 9460 4120 9512
rect 5356 9460 5408 9512
rect 6460 9460 6512 9512
rect 3424 9392 3476 9444
rect 3056 9324 3108 9376
rect 3240 9324 3292 9376
rect 4160 9324 4212 9376
rect 6092 9392 6144 9444
rect 6736 9435 6788 9444
rect 6736 9401 6745 9435
rect 6745 9401 6779 9435
rect 6779 9401 6788 9435
rect 6736 9392 6788 9401
rect 6828 9324 6880 9376
rect 8300 9324 8352 9376
rect 9220 9367 9272 9376
rect 9220 9333 9237 9367
rect 9237 9333 9271 9367
rect 9271 9333 9272 9367
rect 9220 9324 9272 9333
rect 2566 9222 2618 9274
rect 2630 9222 2682 9274
rect 2694 9222 2746 9274
rect 2758 9222 2810 9274
rect 2822 9222 2874 9274
rect 7566 9222 7618 9274
rect 7630 9222 7682 9274
rect 7694 9222 7746 9274
rect 7758 9222 7810 9274
rect 7822 9222 7874 9274
rect 1400 9120 1452 9172
rect 2412 9120 2464 9172
rect 3148 9163 3200 9172
rect 3148 9129 3157 9163
rect 3157 9129 3191 9163
rect 3191 9129 3200 9163
rect 3148 9120 3200 9129
rect 1584 9052 1636 9104
rect 5356 9120 5408 9172
rect 6000 9120 6052 9172
rect 6552 9120 6604 9172
rect 8852 9120 8904 9172
rect 9404 9163 9456 9172
rect 9404 9129 9413 9163
rect 9413 9129 9447 9163
rect 9447 9129 9456 9163
rect 9404 9120 9456 9129
rect 5172 9052 5224 9104
rect 5724 9095 5776 9104
rect 1492 8959 1544 8968
rect 1492 8925 1501 8959
rect 1501 8925 1535 8959
rect 1535 8925 1544 8959
rect 1492 8916 1544 8925
rect 1676 8916 1728 8968
rect 3792 8984 3844 9036
rect 1400 8848 1452 8900
rect 2412 8848 2464 8900
rect 3332 8916 3384 8968
rect 1768 8780 1820 8832
rect 1952 8780 2004 8832
rect 3516 8848 3568 8900
rect 4804 8984 4856 9036
rect 5724 9061 5733 9095
rect 5733 9061 5767 9095
rect 5767 9061 5776 9095
rect 5724 9052 5776 9061
rect 6184 9052 6236 9104
rect 4252 8959 4304 8968
rect 4252 8925 4261 8959
rect 4261 8925 4295 8959
rect 4295 8925 4304 8959
rect 4252 8916 4304 8925
rect 4620 8916 4672 8968
rect 4988 8916 5040 8968
rect 5540 8959 5592 8968
rect 5540 8925 5549 8959
rect 5549 8925 5583 8959
rect 5583 8925 5592 8959
rect 5540 8916 5592 8925
rect 5908 8959 5960 8968
rect 5908 8925 5917 8959
rect 5917 8925 5951 8959
rect 5951 8925 5960 8959
rect 5908 8916 5960 8925
rect 6368 8984 6420 9036
rect 8392 8984 8444 9036
rect 9128 8984 9180 9036
rect 8576 8916 8628 8968
rect 8760 8959 8812 8968
rect 8760 8925 8769 8959
rect 8769 8925 8803 8959
rect 8803 8925 8812 8959
rect 8760 8916 8812 8925
rect 4344 8848 4396 8900
rect 5724 8848 5776 8900
rect 6184 8848 6236 8900
rect 7840 8848 7892 8900
rect 3792 8823 3844 8832
rect 3792 8789 3801 8823
rect 3801 8789 3835 8823
rect 3835 8789 3844 8823
rect 3792 8780 3844 8789
rect 4804 8780 4856 8832
rect 5448 8780 5500 8832
rect 8392 8848 8444 8900
rect 8300 8780 8352 8832
rect 16580 8780 16632 8832
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 5194 8678 5246 8730
rect 5258 8678 5310 8730
rect 5322 8678 5374 8730
rect 3148 8576 3200 8628
rect 3240 8508 3292 8560
rect 1584 8440 1636 8492
rect 1768 8483 1820 8492
rect 1768 8449 1777 8483
rect 1777 8449 1811 8483
rect 1811 8449 1820 8483
rect 1768 8440 1820 8449
rect 3792 8440 3844 8492
rect 5540 8576 5592 8628
rect 4252 8508 4304 8560
rect 1860 8372 1912 8424
rect 2136 8415 2188 8424
rect 2136 8381 2145 8415
rect 2145 8381 2179 8415
rect 2179 8381 2188 8415
rect 2136 8372 2188 8381
rect 4436 8440 4488 8492
rect 4988 8483 5040 8492
rect 4988 8449 4997 8483
rect 4997 8449 5031 8483
rect 5031 8449 5040 8483
rect 4988 8440 5040 8449
rect 5724 8508 5776 8560
rect 6184 8576 6236 8628
rect 8760 8576 8812 8628
rect 9128 8576 9180 8628
rect 7472 8508 7524 8560
rect 5908 8440 5960 8492
rect 6184 8372 6236 8424
rect 6460 8372 6512 8424
rect 8576 8508 8628 8560
rect 16580 8576 16632 8628
rect 8208 8372 8260 8424
rect 8392 8372 8444 8424
rect 8760 8372 8812 8424
rect 4620 8279 4672 8288
rect 4620 8245 4629 8279
rect 4629 8245 4663 8279
rect 4663 8245 4672 8279
rect 4620 8236 4672 8245
rect 5816 8304 5868 8356
rect 6828 8304 6880 8356
rect 5448 8236 5500 8288
rect 6368 8279 6420 8288
rect 6368 8245 6377 8279
rect 6377 8245 6411 8279
rect 6411 8245 6420 8279
rect 6368 8236 6420 8245
rect 7012 8236 7064 8288
rect 7196 8236 7248 8288
rect 9036 8236 9088 8288
rect 2566 8134 2618 8186
rect 2630 8134 2682 8186
rect 2694 8134 2746 8186
rect 2758 8134 2810 8186
rect 2822 8134 2874 8186
rect 7566 8134 7618 8186
rect 7630 8134 7682 8186
rect 7694 8134 7746 8186
rect 7758 8134 7810 8186
rect 7822 8134 7874 8186
rect 2136 8032 2188 8084
rect 4620 8032 4672 8084
rect 9312 8032 9364 8084
rect 2964 7964 3016 8016
rect 3240 7964 3292 8016
rect 2964 7828 3016 7880
rect 7932 7964 7984 8016
rect 8576 7964 8628 8016
rect 5632 7896 5684 7948
rect 6368 7896 6420 7948
rect 7104 7896 7156 7948
rect 4436 7828 4488 7880
rect 5724 7828 5776 7880
rect 7472 7828 7524 7880
rect 8668 7828 8720 7880
rect 8760 7871 8812 7880
rect 8760 7837 8769 7871
rect 8769 7837 8803 7871
rect 8803 7837 8812 7871
rect 8760 7828 8812 7837
rect 6460 7760 6512 7812
rect 3884 7692 3936 7744
rect 7196 7692 7248 7744
rect 7932 7692 7984 7744
rect 8116 7735 8168 7744
rect 8116 7701 8125 7735
rect 8125 7701 8159 7735
rect 8159 7701 8168 7735
rect 8116 7692 8168 7701
rect 8300 7735 8352 7744
rect 8300 7701 8309 7735
rect 8309 7701 8343 7735
rect 8343 7701 8352 7735
rect 8300 7692 8352 7701
rect 8392 7735 8444 7744
rect 8392 7701 8401 7735
rect 8401 7701 8435 7735
rect 8435 7701 8444 7735
rect 8392 7692 8444 7701
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 5194 7590 5246 7642
rect 5258 7590 5310 7642
rect 5322 7590 5374 7642
rect 1400 7531 1452 7540
rect 1400 7497 1409 7531
rect 1409 7497 1443 7531
rect 1443 7497 1452 7531
rect 1400 7488 1452 7497
rect 3424 7488 3476 7540
rect 5632 7488 5684 7540
rect 8392 7488 8444 7540
rect 3148 7420 3200 7472
rect 5448 7420 5500 7472
rect 7472 7420 7524 7472
rect 3884 7395 3936 7404
rect 3884 7361 3893 7395
rect 3893 7361 3927 7395
rect 3927 7361 3936 7395
rect 3884 7352 3936 7361
rect 4804 7352 4856 7404
rect 6828 7352 6880 7404
rect 8208 7395 8260 7404
rect 8208 7361 8217 7395
rect 8217 7361 8251 7395
rect 8251 7361 8260 7395
rect 8208 7352 8260 7361
rect 2412 7284 2464 7336
rect 3056 7284 3108 7336
rect 3424 7327 3476 7336
rect 3424 7293 3433 7327
rect 3433 7293 3467 7327
rect 3467 7293 3476 7327
rect 3424 7284 3476 7293
rect 7012 7284 7064 7336
rect 4804 7216 4856 7268
rect 4988 7216 5040 7268
rect 1676 7191 1728 7200
rect 1676 7157 1685 7191
rect 1685 7157 1719 7191
rect 1719 7157 1728 7191
rect 1676 7148 1728 7157
rect 8300 7148 8352 7200
rect 8944 7148 8996 7200
rect 9036 7191 9088 7200
rect 9036 7157 9045 7191
rect 9045 7157 9079 7191
rect 9079 7157 9088 7191
rect 9036 7148 9088 7157
rect 9312 7148 9364 7200
rect 2566 7046 2618 7098
rect 2630 7046 2682 7098
rect 2694 7046 2746 7098
rect 2758 7046 2810 7098
rect 2822 7046 2874 7098
rect 7566 7046 7618 7098
rect 7630 7046 7682 7098
rect 7694 7046 7746 7098
rect 7758 7046 7810 7098
rect 7822 7046 7874 7098
rect 1676 6944 1728 6996
rect 4436 6944 4488 6996
rect 3424 6808 3476 6860
rect 4160 6876 4212 6928
rect 7196 6876 7248 6928
rect 8116 6876 8168 6928
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 7932 6808 7984 6860
rect 2504 6672 2556 6724
rect 2688 6672 2740 6724
rect 5080 6783 5132 6792
rect 5080 6749 5089 6783
rect 5089 6749 5123 6783
rect 5123 6749 5132 6783
rect 5080 6740 5132 6749
rect 5816 6740 5868 6792
rect 8024 6740 8076 6792
rect 9128 6740 9180 6792
rect 7196 6672 7248 6724
rect 1492 6604 1544 6656
rect 2964 6604 3016 6656
rect 3424 6647 3476 6656
rect 3424 6613 3433 6647
rect 3433 6613 3467 6647
rect 3467 6613 3476 6647
rect 3424 6604 3476 6613
rect 4068 6604 4120 6656
rect 5816 6647 5868 6656
rect 5816 6613 5825 6647
rect 5825 6613 5859 6647
rect 5859 6613 5868 6647
rect 5816 6604 5868 6613
rect 6368 6604 6420 6656
rect 6828 6604 6880 6656
rect 7104 6604 7156 6656
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 5194 6502 5246 6554
rect 5258 6502 5310 6554
rect 5322 6502 5374 6554
rect 1492 6332 1544 6384
rect 2688 6264 2740 6316
rect 3148 6264 3200 6316
rect 3976 6332 4028 6384
rect 5816 6264 5868 6316
rect 6000 6307 6052 6316
rect 6000 6273 6009 6307
rect 6009 6273 6043 6307
rect 6043 6273 6052 6307
rect 6000 6264 6052 6273
rect 6184 6264 6236 6316
rect 7012 6400 7064 6452
rect 7840 6400 7892 6452
rect 6828 6332 6880 6384
rect 7012 6307 7064 6316
rect 1308 6239 1360 6248
rect 1308 6205 1317 6239
rect 1317 6205 1351 6239
rect 1351 6205 1360 6239
rect 1308 6196 1360 6205
rect 3608 6239 3660 6248
rect 3608 6205 3617 6239
rect 3617 6205 3651 6239
rect 3651 6205 3660 6239
rect 3608 6196 3660 6205
rect 5448 6128 5500 6180
rect 7012 6273 7021 6307
rect 7021 6273 7055 6307
rect 7055 6273 7064 6307
rect 7012 6264 7064 6273
rect 7932 6332 7984 6384
rect 8116 6332 8168 6384
rect 6920 6239 6972 6248
rect 6920 6205 6929 6239
rect 6929 6205 6963 6239
rect 6963 6205 6972 6239
rect 6920 6196 6972 6205
rect 9404 6264 9456 6316
rect 8116 6196 8168 6248
rect 8208 6196 8260 6248
rect 7288 6128 7340 6180
rect 1952 6060 2004 6112
rect 4988 6060 5040 6112
rect 6828 6060 6880 6112
rect 9128 6103 9180 6112
rect 9128 6069 9137 6103
rect 9137 6069 9171 6103
rect 9171 6069 9180 6103
rect 9128 6060 9180 6069
rect 2566 5958 2618 6010
rect 2630 5958 2682 6010
rect 2694 5958 2746 6010
rect 2758 5958 2810 6010
rect 2822 5958 2874 6010
rect 7566 5958 7618 6010
rect 7630 5958 7682 6010
rect 7694 5958 7746 6010
rect 7758 5958 7810 6010
rect 7822 5958 7874 6010
rect 1308 5788 1360 5840
rect 4344 5856 4396 5908
rect 5448 5856 5500 5908
rect 6920 5899 6972 5908
rect 4620 5788 4672 5840
rect 6920 5865 6929 5899
rect 6929 5865 6963 5899
rect 6963 5865 6972 5899
rect 6920 5856 6972 5865
rect 7012 5856 7064 5908
rect 8116 5856 8168 5908
rect 8944 5856 8996 5908
rect 11520 5856 11572 5908
rect 9496 5788 9548 5840
rect 3424 5720 3476 5772
rect 3884 5652 3936 5704
rect 6736 5720 6788 5772
rect 1952 5584 2004 5636
rect 3148 5584 3200 5636
rect 3976 5584 4028 5636
rect 6552 5652 6604 5704
rect 4804 5584 4856 5636
rect 5724 5584 5776 5636
rect 6092 5584 6144 5636
rect 7932 5652 7984 5704
rect 8852 5720 8904 5772
rect 8300 5695 8352 5704
rect 8300 5661 8309 5695
rect 8309 5661 8343 5695
rect 8343 5661 8352 5695
rect 8300 5652 8352 5661
rect 9036 5695 9088 5704
rect 8208 5584 8260 5636
rect 9036 5661 9045 5695
rect 9045 5661 9079 5695
rect 9079 5661 9088 5695
rect 9036 5652 9088 5661
rect 8760 5584 8812 5636
rect 3332 5559 3384 5568
rect 3332 5525 3341 5559
rect 3341 5525 3375 5559
rect 3375 5525 3384 5559
rect 3332 5516 3384 5525
rect 6552 5516 6604 5568
rect 7288 5516 7340 5568
rect 7932 5516 7984 5568
rect 8300 5516 8352 5568
rect 8576 5516 8628 5568
rect 9220 5516 9272 5568
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 5194 5414 5246 5466
rect 5258 5414 5310 5466
rect 5322 5414 5374 5466
rect 3608 5312 3660 5364
rect 5724 5355 5776 5364
rect 5724 5321 5733 5355
rect 5733 5321 5767 5355
rect 5767 5321 5776 5355
rect 5724 5312 5776 5321
rect 5908 5312 5960 5364
rect 6736 5312 6788 5364
rect 6276 5244 6328 5296
rect 7380 5244 7432 5296
rect 7656 5312 7708 5364
rect 8852 5287 8904 5296
rect 8852 5253 8861 5287
rect 8861 5253 8895 5287
rect 8895 5253 8904 5287
rect 8852 5244 8904 5253
rect 3424 5219 3476 5228
rect 3424 5185 3433 5219
rect 3433 5185 3467 5219
rect 3467 5185 3476 5219
rect 3424 5176 3476 5185
rect 6644 5176 6696 5228
rect 7932 5219 7984 5228
rect 7932 5185 7941 5219
rect 7941 5185 7975 5219
rect 7975 5185 7984 5219
rect 7932 5176 7984 5185
rect 7288 5108 7340 5160
rect 8392 5176 8444 5228
rect 8576 5176 8628 5228
rect 9220 5219 9272 5228
rect 9220 5185 9229 5219
rect 9229 5185 9263 5219
rect 9263 5185 9272 5219
rect 9220 5176 9272 5185
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 9404 5108 9456 5160
rect 4160 5040 4212 5092
rect 8944 5040 8996 5092
rect 3700 4972 3752 5024
rect 4528 4972 4580 5024
rect 5356 4972 5408 5024
rect 6000 4972 6052 5024
rect 6920 4972 6972 5024
rect 7932 4972 7984 5024
rect 7566 4870 7618 4922
rect 7630 4870 7682 4922
rect 7694 4870 7746 4922
rect 7758 4870 7810 4922
rect 7822 4870 7874 4922
rect 3424 4811 3476 4820
rect 3424 4777 3433 4811
rect 3433 4777 3467 4811
rect 3467 4777 3476 4811
rect 3424 4768 3476 4777
rect 3240 4700 3292 4752
rect 8668 4768 8720 4820
rect 4068 4700 4120 4752
rect 4804 4700 4856 4752
rect 3332 4564 3384 4616
rect 3976 4564 4028 4616
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 5356 4607 5408 4616
rect 5356 4573 5365 4607
rect 5365 4573 5399 4607
rect 5399 4573 5408 4607
rect 5356 4564 5408 4573
rect 7104 4632 7156 4684
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 9128 4564 9180 4616
rect 9404 4607 9456 4616
rect 9404 4573 9413 4607
rect 9413 4573 9447 4607
rect 9447 4573 9456 4607
rect 9404 4564 9456 4573
rect 4436 4496 4488 4548
rect 6092 4496 6144 4548
rect 8116 4496 8168 4548
rect 9220 4496 9272 4548
rect 4252 4471 4304 4480
rect 4252 4437 4261 4471
rect 4261 4437 4295 4471
rect 4295 4437 4304 4471
rect 4252 4428 4304 4437
rect 4344 4428 4396 4480
rect 4988 4428 5040 4480
rect 6644 4428 6696 4480
rect 8668 4428 8720 4480
rect 16580 4428 16632 4480
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 5194 4326 5246 4378
rect 5258 4326 5310 4378
rect 5322 4326 5374 4378
rect 3240 4224 3292 4276
rect 5724 4224 5776 4276
rect 5816 4224 5868 4276
rect 3148 4088 3200 4140
rect 3424 4088 3476 4140
rect 3700 4088 3752 4140
rect 4068 4156 4120 4208
rect 4436 4156 4488 4208
rect 5172 4156 5224 4208
rect 8300 4224 8352 4276
rect 9496 4224 9548 4276
rect 6276 4131 6328 4140
rect 3608 4020 3660 4072
rect 3516 3952 3568 4004
rect 4804 4063 4856 4072
rect 4804 4029 4813 4063
rect 4813 4029 4847 4063
rect 4847 4029 4856 4063
rect 4804 4020 4856 4029
rect 6276 4097 6285 4131
rect 6285 4097 6319 4131
rect 6319 4097 6328 4131
rect 6276 4088 6328 4097
rect 7196 4088 7248 4140
rect 5172 4020 5224 4072
rect 6460 4020 6512 4072
rect 5908 3952 5960 4004
rect 8024 4156 8076 4208
rect 8576 4156 8628 4208
rect 7932 4088 7984 4140
rect 8208 4088 8260 4140
rect 8668 4131 8720 4140
rect 8668 4097 8677 4131
rect 8677 4097 8711 4131
rect 8711 4097 8720 4131
rect 8668 4088 8720 4097
rect 8944 4131 8996 4140
rect 8944 4097 8953 4131
rect 8953 4097 8987 4131
rect 8987 4097 8996 4131
rect 8944 4088 8996 4097
rect 8208 3952 8260 4004
rect 3884 3884 3936 3936
rect 6736 3884 6788 3936
rect 6828 3927 6880 3936
rect 6828 3893 6845 3927
rect 6845 3893 6879 3927
rect 6879 3893 6880 3927
rect 7196 3927 7248 3936
rect 6828 3884 6880 3893
rect 7196 3893 7205 3927
rect 7205 3893 7239 3927
rect 7239 3893 7248 3927
rect 7196 3884 7248 3893
rect 7932 3927 7984 3936
rect 7932 3893 7941 3927
rect 7941 3893 7975 3927
rect 7975 3893 7984 3927
rect 7932 3884 7984 3893
rect 8116 3884 8168 3936
rect 7566 3782 7618 3834
rect 7630 3782 7682 3834
rect 7694 3782 7746 3834
rect 7758 3782 7810 3834
rect 7822 3782 7874 3834
rect 3608 3723 3660 3732
rect 3608 3689 3617 3723
rect 3617 3689 3651 3723
rect 3651 3689 3660 3723
rect 3608 3680 3660 3689
rect 5172 3680 5224 3732
rect 6368 3680 6420 3732
rect 6644 3680 6696 3732
rect 6736 3680 6788 3732
rect 3424 3612 3476 3664
rect 4620 3612 4672 3664
rect 5540 3612 5592 3664
rect 3424 3519 3476 3528
rect 3424 3485 3433 3519
rect 3433 3485 3467 3519
rect 3467 3485 3476 3519
rect 3424 3476 3476 3485
rect 4160 3476 4212 3528
rect 4252 3519 4304 3528
rect 4252 3485 4261 3519
rect 4261 3485 4295 3519
rect 4295 3485 4304 3519
rect 5172 3544 5224 3596
rect 4252 3476 4304 3485
rect 4896 3476 4948 3528
rect 7196 3544 7248 3596
rect 6000 3476 6052 3528
rect 6736 3519 6788 3528
rect 5080 3451 5132 3460
rect 5080 3417 5089 3451
rect 5089 3417 5123 3451
rect 5123 3417 5132 3451
rect 5080 3408 5132 3417
rect 5908 3451 5960 3460
rect 5908 3417 5917 3451
rect 5917 3417 5951 3451
rect 5951 3417 5960 3451
rect 5908 3408 5960 3417
rect 6092 3451 6144 3460
rect 6092 3417 6101 3451
rect 6101 3417 6135 3451
rect 6135 3417 6144 3451
rect 6092 3408 6144 3417
rect 3700 3340 3752 3392
rect 4252 3340 4304 3392
rect 4436 3383 4488 3392
rect 4436 3349 4445 3383
rect 4445 3349 4479 3383
rect 4479 3349 4488 3383
rect 4436 3340 4488 3349
rect 6736 3485 6745 3519
rect 6745 3485 6779 3519
rect 6779 3485 6788 3519
rect 6736 3476 6788 3485
rect 8208 3519 8260 3528
rect 8208 3485 8217 3519
rect 8217 3485 8251 3519
rect 8251 3485 8260 3519
rect 8208 3476 8260 3485
rect 8760 3723 8812 3732
rect 8760 3689 8777 3723
rect 8777 3689 8811 3723
rect 8811 3689 8812 3723
rect 8760 3680 8812 3689
rect 9588 3680 9640 3732
rect 7932 3408 7984 3460
rect 6736 3340 6788 3392
rect 7012 3340 7064 3392
rect 7380 3340 7432 3392
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 5194 3238 5246 3290
rect 5258 3238 5310 3290
rect 5322 3238 5374 3290
rect 3608 3136 3660 3188
rect 3884 3136 3936 3188
rect 4436 3068 4488 3120
rect 3700 3043 3752 3052
rect 3700 3009 3709 3043
rect 3709 3009 3743 3043
rect 3743 3009 3752 3043
rect 3700 3000 3752 3009
rect 5540 3043 5592 3052
rect 4068 2975 4120 2984
rect 4068 2941 4077 2975
rect 4077 2941 4111 2975
rect 4111 2941 4120 2975
rect 4068 2932 4120 2941
rect 5540 3009 5549 3043
rect 5549 3009 5583 3043
rect 5583 3009 5592 3043
rect 5540 3000 5592 3009
rect 6368 3136 6420 3188
rect 7380 3136 7432 3188
rect 6460 3068 6512 3120
rect 7012 3068 7064 3120
rect 8484 3136 8536 3188
rect 8392 3068 8444 3120
rect 9312 3000 9364 3052
rect 9588 3000 9640 3052
rect 4344 2932 4396 2984
rect 3516 2864 3568 2916
rect 4068 2796 4120 2848
rect 6644 2932 6696 2984
rect 8484 2864 8536 2916
rect 6552 2796 6604 2848
rect 9220 2839 9272 2848
rect 9220 2805 9229 2839
rect 9229 2805 9263 2839
rect 9263 2805 9272 2839
rect 9220 2796 9272 2805
rect 7566 2694 7618 2746
rect 7630 2694 7682 2746
rect 7694 2694 7746 2746
rect 7758 2694 7810 2746
rect 7822 2694 7874 2746
rect 4252 2592 4304 2644
rect 4620 2592 4672 2644
rect 5448 2592 5500 2644
rect 6276 2592 6328 2644
rect 8392 2635 8444 2644
rect 8392 2601 8409 2635
rect 8409 2601 8443 2635
rect 8443 2601 8444 2635
rect 8392 2592 8444 2601
rect 3608 2456 3660 2508
rect 4160 2456 4212 2508
rect 3332 2431 3384 2440
rect 3332 2397 3341 2431
rect 3341 2397 3375 2431
rect 3375 2397 3384 2431
rect 3332 2388 3384 2397
rect 7012 2456 7064 2508
rect 5908 2388 5960 2440
rect 6368 2431 6420 2440
rect 6368 2397 6377 2431
rect 6377 2397 6411 2431
rect 6411 2397 6420 2431
rect 6368 2388 6420 2397
rect 8944 2456 8996 2508
rect 9128 2456 9180 2508
rect 4252 2320 4304 2372
rect 6736 2320 6788 2372
rect 9220 2363 9272 2372
rect 9220 2329 9229 2363
rect 9229 2329 9263 2363
rect 9263 2329 9272 2363
rect 9220 2320 9272 2329
rect 9312 2363 9364 2372
rect 9312 2329 9321 2363
rect 9321 2329 9355 2363
rect 9355 2329 9364 2363
rect 9312 2320 9364 2329
rect 9588 2320 9640 2372
rect 4620 2252 4672 2304
rect 5448 2252 5500 2304
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 5194 2150 5246 2202
rect 5258 2150 5310 2202
rect 5322 2150 5374 2202
rect 2688 2048 2740 2100
rect 3792 1980 3844 2032
rect 4528 1980 4580 2032
rect 5540 1980 5592 2032
rect 3332 1912 3384 1964
rect 7288 2048 7340 2100
rect 8668 2048 8720 2100
rect 9036 2091 9088 2100
rect 9036 2057 9045 2091
rect 9045 2057 9079 2091
rect 9079 2057 9088 2091
rect 9036 2048 9088 2057
rect 8484 1912 8536 1964
rect 16580 1912 16632 1964
rect 5448 1844 5500 1896
rect 6460 1844 6512 1896
rect 9404 1887 9456 1896
rect 9404 1853 9413 1887
rect 9413 1853 9447 1887
rect 9447 1853 9456 1887
rect 9404 1844 9456 1853
rect 20628 1776 20680 1828
rect 4896 1708 4948 1760
rect 9220 1751 9272 1760
rect 9220 1717 9229 1751
rect 9229 1717 9263 1751
rect 9263 1717 9272 1751
rect 9220 1708 9272 1717
rect 7566 1606 7618 1658
rect 7630 1606 7682 1658
rect 7694 1606 7746 1658
rect 7758 1606 7810 1658
rect 7822 1606 7874 1658
rect 4620 1504 4672 1556
rect 3332 1411 3384 1420
rect 3332 1377 3341 1411
rect 3341 1377 3375 1411
rect 3375 1377 3384 1411
rect 3332 1368 3384 1377
rect 3976 1368 4028 1420
rect 6368 1504 6420 1556
rect 8668 1504 8720 1556
rect 9312 1504 9364 1556
rect 6736 1436 6788 1488
rect 4988 1300 5040 1352
rect 5448 1300 5500 1352
rect 6460 1300 6512 1352
rect 4252 1232 4304 1284
rect 4896 1232 4948 1284
rect 6644 1232 6696 1284
rect 7012 1164 7064 1216
rect 5066 1062 5118 1114
rect 5130 1062 5182 1114
rect 5194 1062 5246 1114
rect 5258 1062 5310 1114
rect 5322 1062 5374 1114
<< metal2 >>
rect 938 12322 994 13000
rect 1398 12322 1454 13000
rect 1858 12322 1914 13000
rect 938 12294 1348 12322
rect 938 12200 994 12294
rect 1320 11370 1348 12294
rect 1398 12294 1808 12322
rect 1398 12200 1454 12294
rect 1320 11354 1440 11370
rect 1320 11348 1452 11354
rect 1320 11342 1400 11348
rect 1400 11290 1452 11296
rect 1412 9178 1440 11290
rect 1676 11144 1728 11150
rect 1676 11086 1728 11092
rect 1688 10742 1716 11086
rect 1676 10736 1728 10742
rect 1676 10678 1728 10684
rect 1492 10668 1544 10674
rect 1492 10610 1544 10616
rect 1504 10266 1532 10610
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1490 10024 1546 10033
rect 1490 9959 1546 9968
rect 1504 9654 1532 9959
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1400 9172 1452 9178
rect 1400 9114 1452 9120
rect 1504 8974 1532 9590
rect 1584 9104 1636 9110
rect 1584 9046 1636 9052
rect 1492 8968 1544 8974
rect 1492 8910 1544 8916
rect 1400 8900 1452 8906
rect 1400 8842 1452 8848
rect 1412 7546 1440 8842
rect 1596 8498 1624 9046
rect 1688 8974 1716 10678
rect 1676 8968 1728 8974
rect 1676 8910 1728 8916
rect 1780 8922 1808 12294
rect 1858 12294 2176 12322
rect 1858 12200 1914 12294
rect 1860 11552 1912 11558
rect 1860 11494 1912 11500
rect 1872 11286 1900 11494
rect 1860 11280 1912 11286
rect 1860 11222 1912 11228
rect 1872 10606 1900 11222
rect 2148 11014 2176 12294
rect 2318 12200 2374 13000
rect 2778 12200 2834 13000
rect 3238 12200 3294 13000
rect 3698 12200 3754 13000
rect 4158 12322 4214 13000
rect 4080 12294 4214 12322
rect 2332 11286 2360 12200
rect 2792 11626 2820 12200
rect 2780 11620 2832 11626
rect 2780 11562 2832 11568
rect 2566 11452 2874 11472
rect 2566 11450 2572 11452
rect 2628 11450 2652 11452
rect 2708 11450 2732 11452
rect 2788 11450 2812 11452
rect 2868 11450 2874 11452
rect 2628 11398 2630 11450
rect 2810 11398 2812 11450
rect 2566 11396 2572 11398
rect 2628 11396 2652 11398
rect 2708 11396 2732 11398
rect 2788 11396 2812 11398
rect 2868 11396 2874 11398
rect 2566 11376 2874 11396
rect 2412 11348 2464 11354
rect 2412 11290 2464 11296
rect 2320 11280 2372 11286
rect 2320 11222 2372 11228
rect 2424 11150 2452 11290
rect 2964 11280 3016 11286
rect 3252 11234 3280 12200
rect 2964 11222 3016 11228
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 2688 11144 2740 11150
rect 2740 11092 2912 11098
rect 2688 11086 2912 11092
rect 2700 11070 2912 11086
rect 2976 11082 3004 11222
rect 3160 11206 3280 11234
rect 3516 11280 3568 11286
rect 3516 11222 3568 11228
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 2136 11008 2188 11014
rect 2136 10950 2188 10956
rect 2884 10962 2912 11070
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 3068 10962 3096 11018
rect 1964 10674 1992 10950
rect 2884 10934 3096 10962
rect 1952 10668 2004 10674
rect 1952 10610 2004 10616
rect 1860 10600 1912 10606
rect 1860 10542 1912 10548
rect 2136 10600 2188 10606
rect 2136 10542 2188 10548
rect 1872 9722 1900 10542
rect 2148 10198 2176 10542
rect 2566 10364 2874 10384
rect 2566 10362 2572 10364
rect 2628 10362 2652 10364
rect 2708 10362 2732 10364
rect 2788 10362 2812 10364
rect 2868 10362 2874 10364
rect 2628 10310 2630 10362
rect 2810 10310 2812 10362
rect 2566 10308 2572 10310
rect 2628 10308 2652 10310
rect 2708 10308 2732 10310
rect 2788 10308 2812 10310
rect 2868 10308 2874 10310
rect 2566 10288 2874 10308
rect 2136 10192 2188 10198
rect 2136 10134 2188 10140
rect 1860 9716 1912 9722
rect 1860 9658 1912 9664
rect 1872 9058 1900 9658
rect 2566 9276 2874 9296
rect 2566 9274 2572 9276
rect 2628 9274 2652 9276
rect 2708 9274 2732 9276
rect 2788 9274 2812 9276
rect 2868 9274 2874 9276
rect 2628 9222 2630 9274
rect 2810 9222 2812 9274
rect 2566 9220 2572 9222
rect 2628 9220 2652 9222
rect 2708 9220 2732 9222
rect 2788 9220 2812 9222
rect 2868 9220 2874 9222
rect 2566 9200 2874 9220
rect 2412 9172 2464 9178
rect 2412 9114 2464 9120
rect 1872 9030 1992 9058
rect 1780 8894 1900 8922
rect 1768 8832 1820 8838
rect 1768 8774 1820 8780
rect 1780 8498 1808 8774
rect 1584 8492 1636 8498
rect 1584 8434 1636 8440
rect 1768 8492 1820 8498
rect 1768 8434 1820 8440
rect 1872 8430 1900 8894
rect 1964 8838 1992 9030
rect 2424 8906 2452 9114
rect 2412 8900 2464 8906
rect 2412 8842 2464 8848
rect 1952 8832 2004 8838
rect 1952 8774 2004 8780
rect 1860 8424 1912 8430
rect 1860 8366 1912 8372
rect 2136 8424 2188 8430
rect 2136 8366 2188 8372
rect 2148 8090 2176 8366
rect 2566 8188 2874 8208
rect 2566 8186 2572 8188
rect 2628 8186 2652 8188
rect 2708 8186 2732 8188
rect 2788 8186 2812 8188
rect 2868 8186 2874 8188
rect 2628 8134 2630 8186
rect 2810 8134 2812 8186
rect 2566 8132 2572 8134
rect 2628 8132 2652 8134
rect 2708 8132 2732 8134
rect 2788 8132 2812 8134
rect 2868 8132 2874 8134
rect 2566 8112 2874 8132
rect 2136 8084 2188 8090
rect 2136 8026 2188 8032
rect 2976 8022 3004 10934
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 9382 3096 9998
rect 3160 9738 3188 11206
rect 3240 11076 3292 11082
rect 3240 11018 3292 11024
rect 3424 11076 3476 11082
rect 3424 11018 3476 11024
rect 3252 10826 3280 11018
rect 3252 10798 3372 10826
rect 3240 10736 3292 10742
rect 3240 10678 3292 10684
rect 3252 10198 3280 10678
rect 3240 10192 3292 10198
rect 3240 10134 3292 10140
rect 3160 9710 3280 9738
rect 3148 9580 3200 9586
rect 3148 9522 3200 9528
rect 3056 9376 3108 9382
rect 3056 9318 3108 9324
rect 2964 8016 3016 8022
rect 2964 7958 3016 7964
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 1400 7540 1452 7546
rect 1400 7482 1452 7488
rect 2412 7336 2464 7342
rect 2412 7278 2464 7284
rect 1676 7200 1728 7206
rect 1676 7142 1728 7148
rect 1688 7002 1716 7142
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 2424 6914 2452 7278
rect 2566 7100 2874 7120
rect 2566 7098 2572 7100
rect 2628 7098 2652 7100
rect 2708 7098 2732 7100
rect 2788 7098 2812 7100
rect 2868 7098 2874 7100
rect 2628 7046 2630 7098
rect 2810 7046 2812 7098
rect 2566 7044 2572 7046
rect 2628 7044 2652 7046
rect 2708 7044 2732 7046
rect 2788 7044 2812 7046
rect 2868 7044 2874 7046
rect 2566 7024 2874 7044
rect 2424 6886 2544 6914
rect 2516 6730 2544 6886
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2688 6724 2740 6730
rect 2688 6666 2740 6672
rect 1492 6656 1544 6662
rect 1492 6598 1544 6604
rect 1504 6390 1532 6598
rect 1492 6384 1544 6390
rect 1492 6326 1544 6332
rect 2700 6322 2728 6666
rect 2976 6662 3004 7822
rect 3068 7342 3096 9318
rect 3160 9178 3188 9522
rect 3252 9489 3280 9710
rect 3238 9480 3294 9489
rect 3238 9415 3294 9424
rect 3240 9376 3292 9382
rect 3240 9318 3292 9324
rect 3148 9172 3200 9178
rect 3148 9114 3200 9120
rect 3148 8628 3200 8634
rect 3148 8570 3200 8576
rect 3160 7478 3188 8570
rect 3252 8566 3280 9318
rect 3344 8974 3372 10798
rect 3436 9586 3464 11018
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3424 9444 3476 9450
rect 3424 9386 3476 9392
rect 3332 8968 3384 8974
rect 3332 8910 3384 8916
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3240 8016 3292 8022
rect 3240 7958 3292 7964
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3056 7336 3108 7342
rect 3056 7278 3108 7284
rect 2964 6656 3016 6662
rect 2964 6598 3016 6604
rect 2688 6316 2740 6322
rect 2688 6258 2740 6264
rect 3148 6316 3200 6322
rect 3148 6258 3200 6264
rect 1308 6248 1360 6254
rect 1308 6190 1360 6196
rect 1320 5846 1348 6190
rect 1952 6112 2004 6118
rect 1952 6054 2004 6060
rect 1308 5840 1360 5846
rect 1308 5782 1360 5788
rect 1964 5642 1992 6054
rect 2566 6012 2874 6032
rect 2566 6010 2572 6012
rect 2628 6010 2652 6012
rect 2708 6010 2732 6012
rect 2788 6010 2812 6012
rect 2868 6010 2874 6012
rect 2628 5958 2630 6010
rect 2810 5958 2812 6010
rect 2566 5956 2572 5958
rect 2628 5956 2652 5958
rect 2708 5956 2732 5958
rect 2788 5956 2812 5958
rect 2868 5956 2874 5958
rect 2566 5936 2874 5956
rect 3160 5642 3188 6258
rect 1952 5636 2004 5642
rect 1952 5578 2004 5584
rect 3148 5636 3200 5642
rect 3148 5578 3200 5584
rect 3160 4146 3188 5578
rect 3252 4758 3280 7958
rect 3436 7546 3464 9386
rect 3528 8906 3556 11222
rect 3608 11008 3660 11014
rect 3608 10950 3660 10956
rect 3620 10674 3648 10950
rect 3608 10668 3660 10674
rect 3608 10610 3660 10616
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3424 7540 3476 7546
rect 3424 7482 3476 7488
rect 3436 7342 3464 7482
rect 3424 7336 3476 7342
rect 3424 7278 3476 7284
rect 3436 6866 3464 7278
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3436 5778 3464 6598
rect 3608 6248 3660 6254
rect 3608 6190 3660 6196
rect 3424 5772 3476 5778
rect 3424 5714 3476 5720
rect 3332 5568 3384 5574
rect 3332 5510 3384 5516
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3252 4282 3280 4694
rect 3344 4622 3372 5510
rect 3620 5370 3648 6190
rect 3608 5364 3660 5370
rect 3608 5306 3660 5312
rect 3424 5228 3476 5234
rect 3424 5170 3476 5176
rect 3436 4826 3464 5170
rect 3712 5030 3740 12200
rect 3792 10056 3844 10062
rect 3792 9998 3844 10004
rect 3804 9042 3832 9998
rect 4080 9674 4108 12294
rect 4158 12200 4214 12294
rect 4618 12200 4674 13000
rect 5078 12200 5134 13000
rect 5538 12322 5594 13000
rect 5538 12294 5948 12322
rect 5538 12200 5594 12294
rect 4252 11620 4304 11626
rect 4252 11562 4304 11568
rect 4080 9646 4200 9674
rect 4172 9602 4200 9646
rect 3988 9574 4200 9602
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3792 8832 3844 8838
rect 3792 8774 3844 8780
rect 3804 8498 3832 8774
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7410 3924 7686
rect 3884 7404 3936 7410
rect 3884 7346 3936 7352
rect 3988 6474 4016 9574
rect 4068 9512 4120 9518
rect 4068 9454 4120 9460
rect 4080 6662 4108 9454
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4172 6934 4200 9318
rect 4264 9058 4292 11562
rect 4632 11354 4660 12200
rect 4988 11552 5040 11558
rect 4988 11494 5040 11500
rect 4620 11348 4672 11354
rect 4620 11290 4672 11296
rect 4528 11280 4580 11286
rect 4528 11222 4580 11228
rect 4344 11144 4396 11150
rect 4344 11086 4396 11092
rect 4356 10810 4384 11086
rect 4344 10804 4396 10810
rect 4344 10746 4396 10752
rect 4540 9654 4568 11222
rect 4620 11212 4672 11218
rect 4620 11154 4672 11160
rect 4632 10674 4660 11154
rect 4896 11008 4948 11014
rect 4896 10950 4948 10956
rect 4620 10668 4672 10674
rect 4620 10610 4672 10616
rect 4528 9648 4580 9654
rect 4528 9590 4580 9596
rect 4264 9030 4476 9058
rect 4252 8968 4304 8974
rect 4252 8910 4304 8916
rect 4264 8566 4292 8910
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4160 6928 4212 6934
rect 4160 6870 4212 6876
rect 4068 6656 4120 6662
rect 4068 6598 4120 6604
rect 3988 6446 4108 6474
rect 3976 6384 4028 6390
rect 3976 6326 4028 6332
rect 3884 5704 3936 5710
rect 3884 5646 3936 5652
rect 3700 5024 3752 5030
rect 3700 4966 3752 4972
rect 3424 4820 3476 4826
rect 3424 4762 3476 4768
rect 3332 4616 3384 4622
rect 3332 4558 3384 4564
rect 3240 4276 3292 4282
rect 3240 4218 3292 4224
rect 3148 4140 3200 4146
rect 3148 4082 3200 4088
rect 3424 4140 3476 4146
rect 3424 4082 3476 4088
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3436 3670 3464 4082
rect 3608 4072 3660 4078
rect 3608 4014 3660 4020
rect 3712 4026 3740 4082
rect 3516 4004 3568 4010
rect 3516 3946 3568 3952
rect 3424 3664 3476 3670
rect 3424 3606 3476 3612
rect 3424 3528 3476 3534
rect 3422 3496 3424 3505
rect 3476 3496 3478 3505
rect 3422 3431 3478 3440
rect 2686 3360 2742 3369
rect 2686 3295 2742 3304
rect 2700 2106 2728 3295
rect 3528 2922 3556 3946
rect 3620 3738 3648 4014
rect 3712 3998 3832 4026
rect 3608 3732 3660 3738
rect 3608 3674 3660 3680
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3608 3188 3660 3194
rect 3608 3130 3660 3136
rect 3516 2916 3568 2922
rect 3516 2858 3568 2864
rect 3620 2514 3648 3130
rect 3712 3058 3740 3334
rect 3700 3052 3752 3058
rect 3700 2994 3752 3000
rect 3608 2508 3660 2514
rect 3608 2450 3660 2456
rect 3332 2440 3384 2446
rect 3332 2382 3384 2388
rect 2688 2100 2740 2106
rect 2688 2042 2740 2048
rect 3344 1970 3372 2382
rect 3804 2038 3832 3998
rect 3896 3942 3924 5646
rect 3988 5642 4016 6326
rect 3976 5636 4028 5642
rect 3976 5578 4028 5584
rect 4080 4758 4108 6446
rect 4356 5914 4384 8842
rect 4448 8498 4476 9030
rect 4632 8974 4660 10610
rect 4804 10464 4856 10470
rect 4804 10406 4856 10412
rect 4710 9480 4766 9489
rect 4710 9415 4766 9424
rect 4620 8968 4672 8974
rect 4620 8910 4672 8916
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4632 8090 4660 8230
rect 4620 8084 4672 8090
rect 4620 8026 4672 8032
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 4448 7002 4476 7822
rect 4436 6996 4488 7002
rect 4436 6938 4488 6944
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4632 5846 4660 8026
rect 4620 5840 4672 5846
rect 4620 5782 4672 5788
rect 4160 5092 4212 5098
rect 4160 5034 4212 5040
rect 4068 4752 4120 4758
rect 4068 4694 4120 4700
rect 3976 4616 4028 4622
rect 3976 4558 4028 4564
rect 3884 3936 3936 3942
rect 3884 3878 3936 3884
rect 3896 3194 3924 3878
rect 3884 3188 3936 3194
rect 3884 3130 3936 3136
rect 3792 2032 3844 2038
rect 3792 1974 3844 1980
rect 3332 1964 3384 1970
rect 3332 1906 3384 1912
rect 3344 1426 3372 1906
rect 3988 1426 4016 4558
rect 4080 4214 4108 4694
rect 4068 4208 4120 4214
rect 4068 4150 4120 4156
rect 4172 3534 4200 5034
rect 4528 5024 4580 5030
rect 4528 4966 4580 4972
rect 4436 4548 4488 4554
rect 4436 4490 4488 4496
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 4344 4480 4396 4486
rect 4344 4422 4396 4428
rect 4264 3534 4292 4422
rect 4160 3528 4212 3534
rect 4160 3470 4212 3476
rect 4252 3528 4304 3534
rect 4252 3470 4304 3476
rect 4068 2984 4120 2990
rect 4068 2926 4120 2932
rect 4080 2854 4108 2926
rect 4068 2848 4120 2854
rect 4068 2790 4120 2796
rect 4172 2514 4200 3470
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4264 2650 4292 3334
rect 4356 2990 4384 4422
rect 4448 4214 4476 4490
rect 4436 4208 4488 4214
rect 4436 4150 4488 4156
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4448 3126 4476 3334
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4344 2984 4396 2990
rect 4344 2926 4396 2932
rect 4252 2644 4304 2650
rect 4252 2586 4304 2592
rect 4160 2508 4212 2514
rect 4160 2450 4212 2456
rect 4264 2378 4292 2586
rect 4252 2372 4304 2378
rect 4252 2314 4304 2320
rect 3332 1420 3384 1426
rect 3332 1362 3384 1368
rect 3976 1420 4028 1426
rect 3976 1362 4028 1368
rect 4264 1290 4292 2314
rect 4540 2038 4568 4966
rect 4724 4622 4752 9415
rect 4816 9042 4844 10406
rect 4908 10062 4936 10950
rect 4896 10056 4948 10062
rect 4896 9998 4948 10004
rect 4804 9036 4856 9042
rect 4804 8978 4856 8984
rect 5000 8974 5028 11494
rect 5092 11286 5120 12200
rect 5448 11348 5500 11354
rect 5448 11290 5500 11296
rect 5632 11348 5684 11354
rect 5920 11336 5948 12294
rect 5998 12200 6054 13000
rect 6458 12200 6514 13000
rect 9494 12336 9550 12345
rect 9494 12271 9550 12280
rect 6012 11506 6040 12200
rect 6012 11478 6408 11506
rect 5920 11308 6040 11336
rect 5632 11290 5684 11296
rect 5080 11280 5132 11286
rect 5080 11222 5132 11228
rect 5460 11082 5488 11290
rect 5448 11076 5500 11082
rect 5448 11018 5500 11024
rect 5066 10908 5374 10928
rect 5066 10906 5072 10908
rect 5128 10906 5152 10908
rect 5208 10906 5232 10908
rect 5288 10906 5312 10908
rect 5368 10906 5374 10908
rect 5128 10854 5130 10906
rect 5310 10854 5312 10906
rect 5066 10852 5072 10854
rect 5128 10852 5152 10854
rect 5208 10852 5232 10854
rect 5288 10852 5312 10854
rect 5368 10852 5374 10854
rect 5066 10832 5374 10852
rect 5460 10810 5488 11018
rect 5448 10804 5500 10810
rect 5448 10746 5500 10752
rect 5540 10668 5592 10674
rect 5540 10610 5592 10616
rect 5066 9820 5374 9840
rect 5066 9818 5072 9820
rect 5128 9818 5152 9820
rect 5208 9818 5232 9820
rect 5288 9818 5312 9820
rect 5368 9818 5374 9820
rect 5128 9766 5130 9818
rect 5310 9766 5312 9818
rect 5066 9764 5072 9766
rect 5128 9764 5152 9766
rect 5208 9764 5232 9766
rect 5288 9764 5312 9766
rect 5368 9764 5374 9766
rect 5066 9744 5374 9764
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5368 9178 5396 9454
rect 5356 9172 5408 9178
rect 5356 9114 5408 9120
rect 5172 9104 5224 9110
rect 5552 9058 5580 10610
rect 5224 9052 5580 9058
rect 5172 9046 5580 9052
rect 5184 9030 5580 9046
rect 4988 8968 5040 8974
rect 4988 8910 5040 8916
rect 5540 8968 5592 8974
rect 5540 8910 5592 8916
rect 5460 8838 5488 8869
rect 4804 8832 4856 8838
rect 4804 8774 4856 8780
rect 5448 8832 5500 8838
rect 5552 8786 5580 8910
rect 5500 8780 5580 8786
rect 5448 8774 5580 8780
rect 4816 7410 4844 8774
rect 5460 8758 5580 8774
rect 5066 8732 5374 8752
rect 5066 8730 5072 8732
rect 5128 8730 5152 8732
rect 5208 8730 5232 8732
rect 5288 8730 5312 8732
rect 5368 8730 5374 8732
rect 5128 8678 5130 8730
rect 5310 8678 5312 8730
rect 5066 8676 5072 8678
rect 5128 8676 5152 8678
rect 5208 8676 5232 8678
rect 5288 8676 5312 8678
rect 5368 8676 5374 8678
rect 5066 8656 5374 8676
rect 5460 8514 5488 8758
rect 5644 8650 5672 11290
rect 5908 11212 5960 11218
rect 5908 11154 5960 11160
rect 5724 11076 5776 11082
rect 5724 11018 5776 11024
rect 5736 9110 5764 11018
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 9586 5856 10406
rect 5816 9580 5868 9586
rect 5816 9522 5868 9528
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5736 8906 5764 9046
rect 5920 8974 5948 11154
rect 6012 9353 6040 11308
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6184 11144 6236 11150
rect 6184 11086 6236 11092
rect 6104 10742 6132 11086
rect 6196 11014 6224 11086
rect 6184 11008 6236 11014
rect 6184 10950 6236 10956
rect 6092 10736 6144 10742
rect 6092 10678 6144 10684
rect 6104 9450 6132 10678
rect 6196 10674 6224 10950
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6184 10056 6236 10062
rect 6184 9998 6236 10004
rect 6092 9444 6144 9450
rect 6092 9386 6144 9392
rect 5998 9344 6054 9353
rect 5998 9279 6054 9288
rect 6000 9172 6052 9178
rect 6000 9114 6052 9120
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5724 8900 5776 8906
rect 5724 8842 5776 8848
rect 5552 8634 5672 8650
rect 5540 8628 5672 8634
rect 5592 8622 5672 8628
rect 5540 8570 5592 8576
rect 5736 8566 5764 8842
rect 5724 8560 5776 8566
rect 4988 8492 5040 8498
rect 5460 8486 5672 8514
rect 5724 8502 5776 8508
rect 4988 8434 5040 8440
rect 4804 7404 4856 7410
rect 4804 7346 4856 7352
rect 5000 7274 5028 8434
rect 5644 8378 5672 8486
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5644 8350 5764 8378
rect 5448 8288 5500 8294
rect 5448 8230 5500 8236
rect 5066 7644 5374 7664
rect 5066 7642 5072 7644
rect 5128 7642 5152 7644
rect 5208 7642 5232 7644
rect 5288 7642 5312 7644
rect 5368 7642 5374 7644
rect 5128 7590 5130 7642
rect 5310 7590 5312 7642
rect 5066 7588 5072 7590
rect 5128 7588 5152 7590
rect 5208 7588 5232 7590
rect 5288 7588 5312 7590
rect 5368 7588 5374 7590
rect 5066 7568 5374 7588
rect 5460 7562 5488 8230
rect 5632 7948 5684 7954
rect 5632 7890 5684 7896
rect 5460 7534 5580 7562
rect 5644 7546 5672 7890
rect 5736 7886 5764 8350
rect 5816 8356 5868 8362
rect 5816 8298 5868 8304
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5448 7472 5500 7478
rect 5448 7414 5500 7420
rect 4804 7268 4856 7274
rect 4804 7210 4856 7216
rect 4988 7268 5040 7274
rect 4988 7210 5040 7216
rect 4816 5642 4844 7210
rect 5080 6792 5132 6798
rect 5000 6740 5080 6746
rect 5000 6734 5132 6740
rect 5000 6718 5120 6734
rect 5000 6118 5028 6718
rect 5066 6556 5374 6576
rect 5066 6554 5072 6556
rect 5128 6554 5152 6556
rect 5208 6554 5232 6556
rect 5288 6554 5312 6556
rect 5368 6554 5374 6556
rect 5128 6502 5130 6554
rect 5310 6502 5312 6554
rect 5066 6500 5072 6502
rect 5128 6500 5152 6502
rect 5208 6500 5232 6502
rect 5288 6500 5312 6502
rect 5368 6500 5374 6502
rect 5066 6480 5374 6500
rect 5460 6186 5488 7414
rect 5448 6180 5500 6186
rect 5448 6122 5500 6128
rect 4988 6112 5040 6118
rect 4988 6054 5040 6060
rect 5448 5908 5500 5914
rect 5448 5850 5500 5856
rect 4804 5636 4856 5642
rect 4804 5578 4856 5584
rect 4816 4758 4844 5578
rect 5066 5468 5374 5488
rect 5066 5466 5072 5468
rect 5128 5466 5152 5468
rect 5208 5466 5232 5468
rect 5288 5466 5312 5468
rect 5368 5466 5374 5468
rect 5128 5414 5130 5466
rect 5310 5414 5312 5466
rect 5066 5412 5072 5414
rect 5128 5412 5152 5414
rect 5208 5412 5232 5414
rect 5288 5412 5312 5414
rect 5368 5412 5374 5414
rect 5066 5392 5374 5412
rect 5356 5024 5408 5030
rect 5356 4966 5408 4972
rect 4804 4752 4856 4758
rect 4804 4694 4856 4700
rect 5368 4622 5396 4966
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 4724 4321 4752 4558
rect 4988 4480 5040 4486
rect 4988 4422 5040 4428
rect 4710 4312 4766 4321
rect 4710 4247 4766 4256
rect 4804 4072 4856 4078
rect 4804 4014 4856 4020
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4632 2650 4660 3606
rect 4620 2644 4672 2650
rect 4620 2586 4672 2592
rect 4620 2304 4672 2310
rect 4620 2246 4672 2252
rect 4528 2032 4580 2038
rect 4528 1974 4580 1980
rect 4632 1562 4660 2246
rect 4620 1556 4672 1562
rect 4620 1498 4672 1504
rect 4816 1306 4844 4014
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4908 1766 4936 3470
rect 4896 1760 4948 1766
rect 4896 1702 4948 1708
rect 5000 1358 5028 4422
rect 5066 4380 5374 4400
rect 5066 4378 5072 4380
rect 5128 4378 5152 4380
rect 5208 4378 5232 4380
rect 5288 4378 5312 4380
rect 5368 4378 5374 4380
rect 5128 4326 5130 4378
rect 5310 4326 5312 4378
rect 5066 4324 5072 4326
rect 5128 4324 5152 4326
rect 5208 4324 5232 4326
rect 5288 4324 5312 4326
rect 5368 4324 5374 4326
rect 5066 4304 5374 4324
rect 5172 4208 5224 4214
rect 5078 4176 5134 4185
rect 5172 4150 5224 4156
rect 5460 4162 5488 5850
rect 5552 5137 5580 7534
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5736 5642 5764 7822
rect 5828 6798 5856 8298
rect 5816 6792 5868 6798
rect 5816 6734 5868 6740
rect 5816 6656 5868 6662
rect 5816 6598 5868 6604
rect 5828 6322 5856 6598
rect 5816 6316 5868 6322
rect 5816 6258 5868 6264
rect 5724 5636 5776 5642
rect 5724 5578 5776 5584
rect 5920 5370 5948 8434
rect 6012 6322 6040 9114
rect 6196 9110 6224 9998
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6184 9104 6236 9110
rect 6184 9046 6236 9052
rect 6184 8900 6236 8906
rect 6184 8842 6236 8848
rect 6196 8634 6224 8842
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 6196 6322 6224 8366
rect 6288 6866 6316 9522
rect 6380 9160 6408 11478
rect 6472 11234 6500 12200
rect 7566 11452 7874 11472
rect 7566 11450 7572 11452
rect 7628 11450 7652 11452
rect 7708 11450 7732 11452
rect 7788 11450 7812 11452
rect 7868 11450 7874 11452
rect 7628 11398 7630 11450
rect 7810 11398 7812 11450
rect 7566 11396 7572 11398
rect 7628 11396 7652 11398
rect 7708 11396 7732 11398
rect 7788 11396 7812 11398
rect 7868 11396 7874 11398
rect 7566 11376 7874 11396
rect 8116 11348 8168 11354
rect 8116 11290 8168 11296
rect 8668 11348 8720 11354
rect 8668 11290 8720 11296
rect 7932 11280 7984 11286
rect 6472 11206 6684 11234
rect 7932 11222 7984 11228
rect 6460 11144 6512 11150
rect 6460 11086 6512 11092
rect 6472 9518 6500 11086
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6460 9512 6512 9518
rect 6460 9454 6512 9460
rect 6564 9178 6592 9522
rect 6552 9172 6604 9178
rect 6380 9132 6500 9160
rect 6368 9036 6420 9042
rect 6368 8978 6420 8984
rect 6380 8294 6408 8978
rect 6472 8514 6500 9132
rect 6552 9114 6604 9120
rect 6472 8486 6592 8514
rect 6460 8424 6512 8430
rect 6460 8366 6512 8372
rect 6368 8288 6420 8294
rect 6368 8230 6420 8236
rect 6380 7954 6408 8230
rect 6368 7948 6420 7954
rect 6368 7890 6420 7896
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6000 6316 6052 6322
rect 6000 6258 6052 6264
rect 6184 6316 6236 6322
rect 6184 6258 6236 6264
rect 6092 5636 6144 5642
rect 6092 5578 6144 5584
rect 5724 5364 5776 5370
rect 5724 5306 5776 5312
rect 5908 5364 5960 5370
rect 5908 5306 5960 5312
rect 5538 5128 5594 5137
rect 5538 5063 5594 5072
rect 5736 4282 5764 5306
rect 6000 5024 6052 5030
rect 6000 4966 6052 4972
rect 5724 4276 5776 4282
rect 5724 4218 5776 4224
rect 5816 4276 5868 4282
rect 5816 4218 5868 4224
rect 5828 4162 5856 4218
rect 5078 4111 5134 4120
rect 5092 3466 5120 4111
rect 5184 4078 5212 4150
rect 5460 4134 5856 4162
rect 5172 4072 5224 4078
rect 5172 4014 5224 4020
rect 5908 4004 5960 4010
rect 5908 3946 5960 3952
rect 5172 3732 5224 3738
rect 5172 3674 5224 3680
rect 5184 3602 5212 3674
rect 5540 3664 5592 3670
rect 5540 3606 5592 3612
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5080 3460 5132 3466
rect 5080 3402 5132 3408
rect 5066 3292 5374 3312
rect 5066 3290 5072 3292
rect 5128 3290 5152 3292
rect 5208 3290 5232 3292
rect 5288 3290 5312 3292
rect 5368 3290 5374 3292
rect 5128 3238 5130 3290
rect 5310 3238 5312 3290
rect 5066 3236 5072 3238
rect 5128 3236 5152 3238
rect 5208 3236 5232 3238
rect 5288 3236 5312 3238
rect 5368 3236 5374 3238
rect 5066 3216 5374 3236
rect 5552 3058 5580 3606
rect 5920 3466 5948 3946
rect 6012 3534 6040 4966
rect 6104 4554 6132 5578
rect 6288 5302 6316 6802
rect 6380 6662 6408 7890
rect 6472 7818 6500 8366
rect 6460 7812 6512 7818
rect 6460 7754 6512 7760
rect 6368 6656 6420 6662
rect 6368 6598 6420 6604
rect 6564 5710 6592 8486
rect 6552 5704 6604 5710
rect 6552 5646 6604 5652
rect 6564 5574 6592 5646
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6656 5234 6684 11206
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 6920 11076 6972 11082
rect 6920 11018 6972 11024
rect 7012 11076 7064 11082
rect 7012 11018 7064 11024
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6748 10266 6776 10610
rect 6736 10260 6788 10266
rect 6736 10202 6788 10208
rect 6734 10160 6790 10169
rect 6734 10095 6790 10104
rect 6748 9450 6776 10095
rect 6736 9444 6788 9450
rect 6736 9386 6788 9392
rect 6828 9376 6880 9382
rect 6734 9344 6790 9353
rect 6828 9318 6880 9324
rect 6734 9279 6790 9288
rect 6748 5778 6776 9279
rect 6840 8362 6868 9318
rect 6828 8356 6880 8362
rect 6828 8298 6880 8304
rect 6932 7426 6960 11018
rect 7024 9586 7052 11018
rect 7116 10470 7144 11154
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7564 11144 7616 11150
rect 7564 11086 7616 11092
rect 7208 10674 7236 11086
rect 7380 11076 7432 11082
rect 7380 11018 7432 11024
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7104 10464 7156 10470
rect 7104 10406 7156 10412
rect 7288 10464 7340 10470
rect 7288 10406 7340 10412
rect 7012 9580 7064 9586
rect 7012 9522 7064 9528
rect 7012 8288 7064 8294
rect 7012 8230 7064 8236
rect 6840 7410 6960 7426
rect 6828 7404 6960 7410
rect 6880 7398 6960 7404
rect 6828 7346 6880 7352
rect 7024 7342 7052 8230
rect 7116 7954 7144 10406
rect 7196 10260 7248 10266
rect 7196 10202 7248 10208
rect 7208 8294 7236 10202
rect 7300 10130 7328 10406
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7288 9716 7340 9722
rect 7288 9658 7340 9664
rect 7196 8288 7248 8294
rect 7196 8230 7248 8236
rect 7104 7948 7156 7954
rect 7104 7890 7156 7896
rect 7012 7336 7064 7342
rect 7012 7278 7064 7284
rect 7116 6746 7144 7890
rect 7196 7744 7248 7750
rect 7196 7686 7248 7692
rect 7208 6934 7236 7686
rect 7196 6928 7248 6934
rect 7196 6870 7248 6876
rect 7024 6718 7144 6746
rect 7196 6724 7248 6730
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6918 6624 6974 6633
rect 6840 6390 6868 6598
rect 6918 6559 6974 6568
rect 6828 6384 6880 6390
rect 6828 6326 6880 6332
rect 6932 6254 6960 6559
rect 7024 6458 7052 6718
rect 7196 6666 7248 6672
rect 7104 6656 7156 6662
rect 7104 6598 7156 6604
rect 7012 6452 7064 6458
rect 7012 6394 7064 6400
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6920 6248 6972 6254
rect 6920 6190 6972 6196
rect 6828 6112 6880 6118
rect 6828 6054 6880 6060
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 6748 5370 6776 5714
rect 6840 5409 6868 6054
rect 7024 5914 7052 6258
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 7012 5908 7064 5914
rect 7012 5850 7064 5856
rect 6826 5400 6882 5409
rect 6736 5364 6788 5370
rect 6826 5335 6882 5344
rect 6736 5306 6788 5312
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6092 4548 6144 4554
rect 6092 4490 6144 4496
rect 6276 4140 6328 4146
rect 6276 4082 6328 4088
rect 6000 3528 6052 3534
rect 6000 3470 6052 3476
rect 5908 3460 5960 3466
rect 5908 3402 5960 3408
rect 6092 3460 6144 3466
rect 6092 3402 6144 3408
rect 5540 3052 5592 3058
rect 5540 2994 5592 3000
rect 6104 2666 6132 3402
rect 5448 2644 5500 2650
rect 5448 2586 5500 2592
rect 5920 2638 6132 2666
rect 6288 2650 6316 4082
rect 6472 4078 6500 4558
rect 6656 4486 6684 5170
rect 6644 4480 6696 4486
rect 6644 4422 6696 4428
rect 6460 4072 6512 4078
rect 6748 4026 6776 5306
rect 6932 5030 6960 5850
rect 6920 5024 6972 5030
rect 6920 4966 6972 4972
rect 7116 4690 7144 6598
rect 7104 4684 7156 4690
rect 7104 4626 7156 4632
rect 7208 4298 7236 6666
rect 7300 6186 7328 9658
rect 7392 9081 7420 11018
rect 7576 10538 7604 11086
rect 7840 11008 7892 11014
rect 7840 10950 7892 10956
rect 7852 10810 7880 10950
rect 7840 10804 7892 10810
rect 7840 10746 7892 10752
rect 7564 10532 7616 10538
rect 7564 10474 7616 10480
rect 7472 10464 7524 10470
rect 7472 10406 7524 10412
rect 7484 9994 7512 10406
rect 7566 10364 7874 10384
rect 7566 10362 7572 10364
rect 7628 10362 7652 10364
rect 7708 10362 7732 10364
rect 7788 10362 7812 10364
rect 7868 10362 7874 10364
rect 7628 10310 7630 10362
rect 7810 10310 7812 10362
rect 7566 10308 7572 10310
rect 7628 10308 7652 10310
rect 7708 10308 7732 10310
rect 7788 10308 7812 10310
rect 7868 10308 7874 10310
rect 7566 10288 7874 10308
rect 7472 9988 7524 9994
rect 7472 9930 7524 9936
rect 7944 9654 7972 11222
rect 8024 11076 8076 11082
rect 8024 11018 8076 11024
rect 8036 10713 8064 11018
rect 8022 10704 8078 10713
rect 8128 10674 8156 11290
rect 8392 11008 8444 11014
rect 8392 10950 8444 10956
rect 8022 10639 8078 10648
rect 8116 10668 8168 10674
rect 7932 9648 7984 9654
rect 7932 9590 7984 9596
rect 7566 9276 7874 9296
rect 7566 9274 7572 9276
rect 7628 9274 7652 9276
rect 7708 9274 7732 9276
rect 7788 9274 7812 9276
rect 7868 9274 7874 9276
rect 7628 9222 7630 9274
rect 7810 9222 7812 9274
rect 7566 9220 7572 9222
rect 7628 9220 7652 9222
rect 7708 9220 7732 9222
rect 7788 9220 7812 9222
rect 7868 9220 7874 9222
rect 7566 9200 7874 9220
rect 7378 9072 7434 9081
rect 7378 9007 7434 9016
rect 7288 6180 7340 6186
rect 7288 6122 7340 6128
rect 7288 5568 7340 5574
rect 7288 5510 7340 5516
rect 7300 5166 7328 5510
rect 7392 5302 7420 9007
rect 7840 8900 7892 8906
rect 7892 8860 7972 8888
rect 7840 8842 7892 8848
rect 7472 8560 7524 8566
rect 7472 8502 7524 8508
rect 7484 7886 7512 8502
rect 7566 8188 7874 8208
rect 7566 8186 7572 8188
rect 7628 8186 7652 8188
rect 7708 8186 7732 8188
rect 7788 8186 7812 8188
rect 7868 8186 7874 8188
rect 7628 8134 7630 8186
rect 7810 8134 7812 8186
rect 7566 8132 7572 8134
rect 7628 8132 7652 8134
rect 7708 8132 7732 8134
rect 7788 8132 7812 8134
rect 7868 8132 7874 8134
rect 7566 8112 7874 8132
rect 7944 8022 7972 8860
rect 7932 8016 7984 8022
rect 7932 7958 7984 7964
rect 7472 7880 7524 7886
rect 7472 7822 7524 7828
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7484 5386 7512 7414
rect 7566 7100 7874 7120
rect 7566 7098 7572 7100
rect 7628 7098 7652 7100
rect 7708 7098 7732 7100
rect 7788 7098 7812 7100
rect 7868 7098 7874 7100
rect 7628 7046 7630 7098
rect 7810 7046 7812 7098
rect 7566 7044 7572 7046
rect 7628 7044 7652 7046
rect 7708 7044 7732 7046
rect 7788 7044 7812 7046
rect 7868 7044 7874 7046
rect 7566 7024 7874 7044
rect 7944 6866 7972 7686
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7840 6452 7892 6458
rect 7840 6394 7892 6400
rect 7852 6202 7880 6394
rect 7944 6390 7972 6802
rect 8036 6798 8064 10639
rect 8116 10610 8168 10616
rect 8404 10606 8432 10950
rect 8392 10600 8444 10606
rect 8392 10542 8444 10548
rect 8116 10464 8168 10470
rect 8116 10406 8168 10412
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8128 9586 8156 10406
rect 8208 10192 8260 10198
rect 8208 10134 8260 10140
rect 8220 9722 8248 10134
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8312 9382 8340 10406
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8404 9194 8432 10542
rect 8484 10056 8536 10062
rect 8484 9998 8536 10004
rect 8220 9166 8432 9194
rect 8220 8430 8248 9166
rect 8404 9042 8432 9166
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8392 8900 8444 8906
rect 8392 8842 8444 8848
rect 8300 8832 8352 8838
rect 8300 8774 8352 8780
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8312 7750 8340 8774
rect 8404 8430 8432 8842
rect 8392 8424 8444 8430
rect 8392 8366 8444 8372
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8128 7041 8156 7686
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8114 7032 8170 7041
rect 8114 6967 8170 6976
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 8024 6792 8076 6798
rect 8024 6734 8076 6740
rect 8128 6390 8156 6870
rect 7932 6384 7984 6390
rect 7932 6326 7984 6332
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8220 6254 8248 7346
rect 8312 7290 8340 7686
rect 8404 7546 8432 7686
rect 8392 7540 8444 7546
rect 8392 7482 8444 7488
rect 8312 7262 8432 7290
rect 8300 7200 8352 7206
rect 8300 7142 8352 7148
rect 8116 6248 8168 6254
rect 7852 6174 7972 6202
rect 8116 6190 8168 6196
rect 8208 6248 8260 6254
rect 8208 6190 8260 6196
rect 7566 6012 7874 6032
rect 7566 6010 7572 6012
rect 7628 6010 7652 6012
rect 7708 6010 7732 6012
rect 7788 6010 7812 6012
rect 7868 6010 7874 6012
rect 7628 5958 7630 6010
rect 7810 5958 7812 6010
rect 7566 5956 7572 5958
rect 7628 5956 7652 5958
rect 7708 5956 7732 5958
rect 7788 5956 7812 5958
rect 7868 5956 7874 5958
rect 7566 5936 7874 5956
rect 7944 5710 7972 6174
rect 8128 5914 8156 6190
rect 8116 5908 8168 5914
rect 8116 5850 8168 5856
rect 8312 5710 8340 7142
rect 7932 5704 7984 5710
rect 7932 5646 7984 5652
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8208 5636 8260 5642
rect 8208 5578 8260 5584
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 7484 5370 7696 5386
rect 7484 5364 7708 5370
rect 7484 5358 7656 5364
rect 7656 5306 7708 5312
rect 7380 5296 7432 5302
rect 7380 5238 7432 5244
rect 7944 5234 7972 5510
rect 7932 5228 7984 5234
rect 7932 5170 7984 5176
rect 7288 5160 7340 5166
rect 7288 5102 7340 5108
rect 7944 5114 7972 5170
rect 6460 4014 6512 4020
rect 6656 3998 6776 4026
rect 7024 4270 7236 4298
rect 6656 3738 6684 3998
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6828 3936 6880 3942
rect 6828 3878 6880 3884
rect 6748 3738 6776 3878
rect 6368 3732 6420 3738
rect 6368 3674 6420 3680
rect 6644 3732 6696 3738
rect 6644 3674 6696 3680
rect 6736 3732 6788 3738
rect 6736 3674 6788 3680
rect 6380 3194 6408 3674
rect 6736 3528 6788 3534
rect 6736 3470 6788 3476
rect 6748 3398 6776 3470
rect 6736 3392 6788 3398
rect 6840 3369 6868 3878
rect 7024 3398 7052 4270
rect 7196 4140 7248 4146
rect 7196 4082 7248 4088
rect 7208 3942 7236 4082
rect 7196 3936 7248 3942
rect 7196 3878 7248 3884
rect 7208 3602 7236 3878
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7300 3505 7328 5102
rect 7944 5086 8064 5114
rect 7932 5024 7984 5030
rect 7932 4966 7984 4972
rect 7566 4924 7874 4944
rect 7566 4922 7572 4924
rect 7628 4922 7652 4924
rect 7708 4922 7732 4924
rect 7788 4922 7812 4924
rect 7868 4922 7874 4924
rect 7628 4870 7630 4922
rect 7810 4870 7812 4922
rect 7566 4868 7572 4870
rect 7628 4868 7652 4870
rect 7708 4868 7732 4870
rect 7788 4868 7812 4870
rect 7868 4868 7874 4870
rect 7566 4848 7874 4868
rect 7944 4146 7972 4966
rect 8036 4214 8064 5086
rect 8116 4548 8168 4554
rect 8116 4490 8168 4496
rect 8024 4208 8076 4214
rect 8024 4150 8076 4156
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 8128 3942 8156 4490
rect 8220 4146 8248 5578
rect 8300 5568 8352 5574
rect 8300 5510 8352 5516
rect 8312 4706 8340 5510
rect 8404 5234 8432 7262
rect 8392 5228 8444 5234
rect 8392 5170 8444 5176
rect 8312 4678 8432 4706
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 8312 4282 8340 4558
rect 8300 4276 8352 4282
rect 8300 4218 8352 4224
rect 8208 4140 8260 4146
rect 8208 4082 8260 4088
rect 8208 4004 8260 4010
rect 8208 3946 8260 3952
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 8116 3936 8168 3942
rect 8116 3878 8168 3884
rect 7566 3836 7874 3856
rect 7566 3834 7572 3836
rect 7628 3834 7652 3836
rect 7708 3834 7732 3836
rect 7788 3834 7812 3836
rect 7868 3834 7874 3836
rect 7628 3782 7630 3834
rect 7810 3782 7812 3834
rect 7566 3780 7572 3782
rect 7628 3780 7652 3782
rect 7708 3780 7732 3782
rect 7788 3780 7812 3782
rect 7868 3780 7874 3782
rect 7566 3760 7874 3780
rect 7286 3496 7342 3505
rect 7944 3466 7972 3878
rect 8220 3534 8248 3946
rect 8208 3528 8260 3534
rect 8208 3470 8260 3476
rect 7286 3431 7342 3440
rect 7932 3460 7984 3466
rect 7012 3392 7064 3398
rect 6736 3334 6788 3340
rect 6826 3360 6882 3369
rect 7012 3334 7064 3340
rect 6826 3295 6882 3304
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6460 3120 6512 3126
rect 6460 3062 6512 3068
rect 7012 3120 7064 3126
rect 7012 3062 7064 3068
rect 6276 2644 6328 2650
rect 5460 2394 5488 2586
rect 5920 2446 5948 2638
rect 6276 2586 6328 2592
rect 5908 2440 5960 2446
rect 5460 2366 5580 2394
rect 5908 2382 5960 2388
rect 6368 2440 6420 2446
rect 6368 2382 6420 2388
rect 5448 2304 5500 2310
rect 5448 2246 5500 2252
rect 5066 2204 5374 2224
rect 5066 2202 5072 2204
rect 5128 2202 5152 2204
rect 5208 2202 5232 2204
rect 5288 2202 5312 2204
rect 5368 2202 5374 2204
rect 5128 2150 5130 2202
rect 5310 2150 5312 2202
rect 5066 2148 5072 2150
rect 5128 2148 5152 2150
rect 5208 2148 5232 2150
rect 5288 2148 5312 2150
rect 5368 2148 5374 2150
rect 5066 2128 5374 2148
rect 5460 1902 5488 2246
rect 5552 2038 5580 2366
rect 5540 2032 5592 2038
rect 5540 1974 5592 1980
rect 5448 1896 5500 1902
rect 5448 1838 5500 1844
rect 5460 1358 5488 1838
rect 6380 1562 6408 2382
rect 6472 1902 6500 3062
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6552 2848 6604 2854
rect 6552 2790 6604 2796
rect 6564 2553 6592 2790
rect 6550 2544 6606 2553
rect 6550 2479 6606 2488
rect 6460 1896 6512 1902
rect 6460 1838 6512 1844
rect 6368 1556 6420 1562
rect 6368 1498 6420 1504
rect 6472 1358 6500 1838
rect 4988 1352 5040 1358
rect 4816 1290 4936 1306
rect 4988 1294 5040 1300
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 6460 1352 6512 1358
rect 6460 1294 6512 1300
rect 6656 1290 6684 2926
rect 7024 2514 7052 3062
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 6736 2372 6788 2378
rect 6736 2314 6788 2320
rect 6748 1494 6776 2314
rect 6736 1488 6788 1494
rect 6736 1430 6788 1436
rect 4252 1284 4304 1290
rect 4816 1284 4948 1290
rect 4816 1278 4896 1284
rect 4252 1226 4304 1232
rect 4896 1226 4948 1232
rect 6644 1284 6696 1290
rect 6644 1226 6696 1232
rect 7024 1222 7052 2450
rect 7300 2106 7328 3431
rect 7932 3402 7984 3408
rect 7380 3392 7432 3398
rect 7380 3334 7432 3340
rect 7392 3194 7420 3334
rect 7380 3188 7432 3194
rect 7380 3130 7432 3136
rect 8404 3126 8432 4678
rect 8496 3194 8524 9998
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8588 8566 8616 8910
rect 8576 8560 8628 8566
rect 8576 8502 8628 8508
rect 8576 8016 8628 8022
rect 8576 7958 8628 7964
rect 8588 5574 8616 7958
rect 8680 7886 8708 11290
rect 9312 10668 9364 10674
rect 9312 10610 9364 10616
rect 9220 9376 9272 9382
rect 9220 9318 9272 9324
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8772 8634 8800 8910
rect 8760 8628 8812 8634
rect 8760 8570 8812 8576
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8772 7886 8800 8366
rect 8668 7880 8720 7886
rect 8668 7822 8720 7828
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8864 5930 8892 9114
rect 9128 9036 9180 9042
rect 9128 8978 9180 8984
rect 9140 8634 9168 8978
rect 9128 8628 9180 8634
rect 9128 8570 9180 8576
rect 9036 8288 9088 8294
rect 9140 8265 9168 8570
rect 9036 8230 9088 8236
rect 9126 8256 9182 8265
rect 9048 7206 9076 8230
rect 9126 8191 9182 8200
rect 9232 7857 9260 9318
rect 9324 8090 9352 10610
rect 9508 10130 9536 12271
rect 16578 11928 16634 11937
rect 16578 11863 16634 11872
rect 16592 11286 16620 11863
rect 20718 11520 20774 11529
rect 20718 11455 20774 11464
rect 16580 11280 16632 11286
rect 16580 11222 16632 11228
rect 16578 11112 16634 11121
rect 16578 11047 16634 11056
rect 16592 10470 16620 11047
rect 16580 10464 16632 10470
rect 16580 10406 16632 10412
rect 9496 10124 9548 10130
rect 9496 10066 9548 10072
rect 9404 10056 9456 10062
rect 9404 9998 9456 10004
rect 9416 9178 9444 9998
rect 9508 9722 9536 10066
rect 9496 9716 9548 9722
rect 9496 9658 9548 9664
rect 16672 9716 16724 9722
rect 16672 9658 16724 9664
rect 16578 9480 16634 9489
rect 16578 9415 16634 9424
rect 9404 9172 9456 9178
rect 9404 9114 9456 9120
rect 16592 8838 16620 9415
rect 16580 8832 16632 8838
rect 16580 8774 16632 8780
rect 16578 8664 16634 8673
rect 16578 8599 16580 8608
rect 16632 8599 16634 8608
rect 16580 8570 16632 8576
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9218 7848 9274 7857
rect 9218 7783 9274 7792
rect 16684 7449 16712 9658
rect 16670 7440 16726 7449
rect 16670 7375 16726 7384
rect 8944 7200 8996 7206
rect 8944 7142 8996 7148
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9312 7200 9364 7206
rect 9312 7142 9364 7148
rect 8680 5902 8892 5930
rect 8956 5914 8984 7142
rect 9048 6882 9076 7142
rect 9048 6854 9260 6882
rect 9128 6792 9180 6798
rect 9128 6734 9180 6740
rect 9140 6118 9168 6734
rect 9232 6225 9260 6854
rect 9218 6216 9274 6225
rect 9218 6151 9274 6160
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 8944 5908 8996 5914
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8588 4214 8616 5170
rect 8680 4826 8708 5902
rect 8944 5850 8996 5856
rect 8852 5772 8904 5778
rect 8852 5714 8904 5720
rect 8760 5636 8812 5642
rect 8760 5578 8812 5584
rect 8668 4820 8720 4826
rect 8668 4762 8720 4768
rect 8772 4593 8800 5578
rect 8864 5302 8892 5714
rect 9036 5704 9088 5710
rect 9036 5646 9088 5652
rect 8852 5296 8904 5302
rect 8852 5238 8904 5244
rect 8944 5092 8996 5098
rect 8944 5034 8996 5040
rect 8758 4584 8814 4593
rect 8758 4519 8814 4528
rect 8668 4480 8720 4486
rect 8668 4422 8720 4428
rect 8576 4208 8628 4214
rect 8576 4150 8628 4156
rect 8680 4146 8708 4422
rect 8668 4140 8720 4146
rect 8668 4082 8720 4088
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8392 3120 8444 3126
rect 8392 3062 8444 3068
rect 8390 2952 8446 2961
rect 8390 2887 8446 2896
rect 8484 2916 8536 2922
rect 7566 2748 7874 2768
rect 7566 2746 7572 2748
rect 7628 2746 7652 2748
rect 7708 2746 7732 2748
rect 7788 2746 7812 2748
rect 7868 2746 7874 2748
rect 7628 2694 7630 2746
rect 7810 2694 7812 2746
rect 7566 2692 7572 2694
rect 7628 2692 7652 2694
rect 7708 2692 7732 2694
rect 7788 2692 7812 2694
rect 7868 2692 7874 2694
rect 7566 2672 7874 2692
rect 8404 2650 8432 2887
rect 8484 2858 8536 2864
rect 8392 2644 8444 2650
rect 8392 2586 8444 2592
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 8496 1970 8524 2858
rect 8680 2106 8708 4082
rect 8772 3738 8800 4519
rect 8956 4146 8984 5034
rect 8944 4140 8996 4146
rect 8944 4082 8996 4088
rect 8760 3732 8812 3738
rect 8760 3674 8812 3680
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 8956 2514 8984 3334
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 9048 2106 9076 5646
rect 9140 4622 9168 6054
rect 9232 5574 9260 6151
rect 9220 5568 9272 5574
rect 9220 5510 9272 5516
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9128 4616 9180 4622
rect 9128 4558 9180 4564
rect 9232 4554 9260 5170
rect 9220 4548 9272 4554
rect 9220 4490 9272 4496
rect 9324 3058 9352 7142
rect 9404 6316 9456 6322
rect 9404 6258 9456 6264
rect 9416 5166 9444 6258
rect 11520 5908 11572 5914
rect 11520 5850 11572 5856
rect 9496 5840 9548 5846
rect 9496 5782 9548 5788
rect 9586 5808 9642 5817
rect 9508 5234 9536 5782
rect 9586 5743 9642 5752
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9404 5160 9456 5166
rect 9404 5102 9456 5108
rect 9404 4616 9456 4622
rect 9404 4558 9456 4564
rect 9312 3052 9364 3058
rect 9312 2994 9364 3000
rect 9220 2848 9272 2854
rect 9220 2790 9272 2796
rect 9128 2508 9180 2514
rect 9128 2450 9180 2456
rect 8668 2100 8720 2106
rect 8668 2042 8720 2048
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 8484 1964 8536 1970
rect 8484 1906 8536 1912
rect 7566 1660 7874 1680
rect 7566 1658 7572 1660
rect 7628 1658 7652 1660
rect 7708 1658 7732 1660
rect 7788 1658 7812 1660
rect 7868 1658 7874 1660
rect 7628 1606 7630 1658
rect 7810 1606 7812 1658
rect 7566 1604 7572 1606
rect 7628 1604 7652 1606
rect 7708 1604 7732 1606
rect 7788 1604 7812 1606
rect 7868 1604 7874 1606
rect 7566 1584 7874 1604
rect 8680 1562 8708 2042
rect 8668 1556 8720 1562
rect 8668 1498 8720 1504
rect 7012 1216 7064 1222
rect 7012 1158 7064 1164
rect 5066 1116 5374 1136
rect 5066 1114 5072 1116
rect 5128 1114 5152 1116
rect 5208 1114 5232 1116
rect 5288 1114 5312 1116
rect 5368 1114 5374 1116
rect 5128 1062 5130 1114
rect 5310 1062 5312 1114
rect 5066 1060 5072 1062
rect 5128 1060 5152 1062
rect 5208 1060 5232 1062
rect 5288 1060 5312 1062
rect 5368 1060 5374 1062
rect 5066 1040 5374 1060
rect 9140 921 9168 2450
rect 9232 2378 9260 2790
rect 9220 2372 9272 2378
rect 9220 2314 9272 2320
rect 9312 2372 9364 2378
rect 9312 2314 9364 2320
rect 9220 1760 9272 1766
rect 9220 1702 9272 1708
rect 9126 912 9182 921
rect 9126 847 9182 856
rect 9232 513 9260 1702
rect 9324 1562 9352 2314
rect 9416 1902 9444 4558
rect 9496 4276 9548 4282
rect 9496 4218 9548 4224
rect 9404 1896 9456 1902
rect 9404 1838 9456 1844
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9416 1329 9444 1838
rect 9508 1737 9536 4218
rect 9600 3738 9628 5743
rect 11532 3777 11560 5850
rect 16580 4480 16632 4486
rect 16580 4422 16632 4428
rect 16592 4185 16620 4422
rect 16578 4176 16634 4185
rect 20732 4162 20760 11455
rect 16578 4111 16634 4120
rect 20640 4134 20760 4162
rect 11518 3768 11574 3777
rect 9588 3732 9640 3738
rect 11518 3703 11574 3712
rect 9588 3674 9640 3680
rect 9600 3058 9628 3674
rect 9588 3052 9640 3058
rect 9588 2994 9640 3000
rect 9600 2378 9628 2994
rect 9588 2372 9640 2378
rect 9588 2314 9640 2320
rect 16578 2136 16634 2145
rect 16578 2071 16634 2080
rect 16592 1970 16620 2071
rect 16580 1964 16632 1970
rect 16580 1906 16632 1912
rect 20640 1834 20668 4134
rect 20628 1828 20680 1834
rect 20628 1770 20680 1776
rect 9494 1728 9550 1737
rect 9494 1663 9550 1672
rect 9402 1320 9458 1329
rect 9402 1255 9458 1264
rect 9218 504 9274 513
rect 9218 439 9274 448
<< via2 >>
rect 1490 9968 1546 10024
rect 2572 11450 2628 11452
rect 2652 11450 2708 11452
rect 2732 11450 2788 11452
rect 2812 11450 2868 11452
rect 2572 11398 2618 11450
rect 2618 11398 2628 11450
rect 2652 11398 2682 11450
rect 2682 11398 2694 11450
rect 2694 11398 2708 11450
rect 2732 11398 2746 11450
rect 2746 11398 2758 11450
rect 2758 11398 2788 11450
rect 2812 11398 2822 11450
rect 2822 11398 2868 11450
rect 2572 11396 2628 11398
rect 2652 11396 2708 11398
rect 2732 11396 2788 11398
rect 2812 11396 2868 11398
rect 2572 10362 2628 10364
rect 2652 10362 2708 10364
rect 2732 10362 2788 10364
rect 2812 10362 2868 10364
rect 2572 10310 2618 10362
rect 2618 10310 2628 10362
rect 2652 10310 2682 10362
rect 2682 10310 2694 10362
rect 2694 10310 2708 10362
rect 2732 10310 2746 10362
rect 2746 10310 2758 10362
rect 2758 10310 2788 10362
rect 2812 10310 2822 10362
rect 2822 10310 2868 10362
rect 2572 10308 2628 10310
rect 2652 10308 2708 10310
rect 2732 10308 2788 10310
rect 2812 10308 2868 10310
rect 2572 9274 2628 9276
rect 2652 9274 2708 9276
rect 2732 9274 2788 9276
rect 2812 9274 2868 9276
rect 2572 9222 2618 9274
rect 2618 9222 2628 9274
rect 2652 9222 2682 9274
rect 2682 9222 2694 9274
rect 2694 9222 2708 9274
rect 2732 9222 2746 9274
rect 2746 9222 2758 9274
rect 2758 9222 2788 9274
rect 2812 9222 2822 9274
rect 2822 9222 2868 9274
rect 2572 9220 2628 9222
rect 2652 9220 2708 9222
rect 2732 9220 2788 9222
rect 2812 9220 2868 9222
rect 2572 8186 2628 8188
rect 2652 8186 2708 8188
rect 2732 8186 2788 8188
rect 2812 8186 2868 8188
rect 2572 8134 2618 8186
rect 2618 8134 2628 8186
rect 2652 8134 2682 8186
rect 2682 8134 2694 8186
rect 2694 8134 2708 8186
rect 2732 8134 2746 8186
rect 2746 8134 2758 8186
rect 2758 8134 2788 8186
rect 2812 8134 2822 8186
rect 2822 8134 2868 8186
rect 2572 8132 2628 8134
rect 2652 8132 2708 8134
rect 2732 8132 2788 8134
rect 2812 8132 2868 8134
rect 2572 7098 2628 7100
rect 2652 7098 2708 7100
rect 2732 7098 2788 7100
rect 2812 7098 2868 7100
rect 2572 7046 2618 7098
rect 2618 7046 2628 7098
rect 2652 7046 2682 7098
rect 2682 7046 2694 7098
rect 2694 7046 2708 7098
rect 2732 7046 2746 7098
rect 2746 7046 2758 7098
rect 2758 7046 2788 7098
rect 2812 7046 2822 7098
rect 2822 7046 2868 7098
rect 2572 7044 2628 7046
rect 2652 7044 2708 7046
rect 2732 7044 2788 7046
rect 2812 7044 2868 7046
rect 3238 9424 3294 9480
rect 2572 6010 2628 6012
rect 2652 6010 2708 6012
rect 2732 6010 2788 6012
rect 2812 6010 2868 6012
rect 2572 5958 2618 6010
rect 2618 5958 2628 6010
rect 2652 5958 2682 6010
rect 2682 5958 2694 6010
rect 2694 5958 2708 6010
rect 2732 5958 2746 6010
rect 2746 5958 2758 6010
rect 2758 5958 2788 6010
rect 2812 5958 2822 6010
rect 2822 5958 2868 6010
rect 2572 5956 2628 5958
rect 2652 5956 2708 5958
rect 2732 5956 2788 5958
rect 2812 5956 2868 5958
rect 3422 3476 3424 3496
rect 3424 3476 3476 3496
rect 3476 3476 3478 3496
rect 3422 3440 3478 3476
rect 2686 3304 2742 3360
rect 4710 9424 4766 9480
rect 9494 12280 9550 12336
rect 5072 10906 5128 10908
rect 5152 10906 5208 10908
rect 5232 10906 5288 10908
rect 5312 10906 5368 10908
rect 5072 10854 5118 10906
rect 5118 10854 5128 10906
rect 5152 10854 5182 10906
rect 5182 10854 5194 10906
rect 5194 10854 5208 10906
rect 5232 10854 5246 10906
rect 5246 10854 5258 10906
rect 5258 10854 5288 10906
rect 5312 10854 5322 10906
rect 5322 10854 5368 10906
rect 5072 10852 5128 10854
rect 5152 10852 5208 10854
rect 5232 10852 5288 10854
rect 5312 10852 5368 10854
rect 5072 9818 5128 9820
rect 5152 9818 5208 9820
rect 5232 9818 5288 9820
rect 5312 9818 5368 9820
rect 5072 9766 5118 9818
rect 5118 9766 5128 9818
rect 5152 9766 5182 9818
rect 5182 9766 5194 9818
rect 5194 9766 5208 9818
rect 5232 9766 5246 9818
rect 5246 9766 5258 9818
rect 5258 9766 5288 9818
rect 5312 9766 5322 9818
rect 5322 9766 5368 9818
rect 5072 9764 5128 9766
rect 5152 9764 5208 9766
rect 5232 9764 5288 9766
rect 5312 9764 5368 9766
rect 5072 8730 5128 8732
rect 5152 8730 5208 8732
rect 5232 8730 5288 8732
rect 5312 8730 5368 8732
rect 5072 8678 5118 8730
rect 5118 8678 5128 8730
rect 5152 8678 5182 8730
rect 5182 8678 5194 8730
rect 5194 8678 5208 8730
rect 5232 8678 5246 8730
rect 5246 8678 5258 8730
rect 5258 8678 5288 8730
rect 5312 8678 5322 8730
rect 5322 8678 5368 8730
rect 5072 8676 5128 8678
rect 5152 8676 5208 8678
rect 5232 8676 5288 8678
rect 5312 8676 5368 8678
rect 5998 9288 6054 9344
rect 5072 7642 5128 7644
rect 5152 7642 5208 7644
rect 5232 7642 5288 7644
rect 5312 7642 5368 7644
rect 5072 7590 5118 7642
rect 5118 7590 5128 7642
rect 5152 7590 5182 7642
rect 5182 7590 5194 7642
rect 5194 7590 5208 7642
rect 5232 7590 5246 7642
rect 5246 7590 5258 7642
rect 5258 7590 5288 7642
rect 5312 7590 5322 7642
rect 5322 7590 5368 7642
rect 5072 7588 5128 7590
rect 5152 7588 5208 7590
rect 5232 7588 5288 7590
rect 5312 7588 5368 7590
rect 5072 6554 5128 6556
rect 5152 6554 5208 6556
rect 5232 6554 5288 6556
rect 5312 6554 5368 6556
rect 5072 6502 5118 6554
rect 5118 6502 5128 6554
rect 5152 6502 5182 6554
rect 5182 6502 5194 6554
rect 5194 6502 5208 6554
rect 5232 6502 5246 6554
rect 5246 6502 5258 6554
rect 5258 6502 5288 6554
rect 5312 6502 5322 6554
rect 5322 6502 5368 6554
rect 5072 6500 5128 6502
rect 5152 6500 5208 6502
rect 5232 6500 5288 6502
rect 5312 6500 5368 6502
rect 5072 5466 5128 5468
rect 5152 5466 5208 5468
rect 5232 5466 5288 5468
rect 5312 5466 5368 5468
rect 5072 5414 5118 5466
rect 5118 5414 5128 5466
rect 5152 5414 5182 5466
rect 5182 5414 5194 5466
rect 5194 5414 5208 5466
rect 5232 5414 5246 5466
rect 5246 5414 5258 5466
rect 5258 5414 5288 5466
rect 5312 5414 5322 5466
rect 5322 5414 5368 5466
rect 5072 5412 5128 5414
rect 5152 5412 5208 5414
rect 5232 5412 5288 5414
rect 5312 5412 5368 5414
rect 4710 4256 4766 4312
rect 5072 4378 5128 4380
rect 5152 4378 5208 4380
rect 5232 4378 5288 4380
rect 5312 4378 5368 4380
rect 5072 4326 5118 4378
rect 5118 4326 5128 4378
rect 5152 4326 5182 4378
rect 5182 4326 5194 4378
rect 5194 4326 5208 4378
rect 5232 4326 5246 4378
rect 5246 4326 5258 4378
rect 5258 4326 5288 4378
rect 5312 4326 5322 4378
rect 5322 4326 5368 4378
rect 5072 4324 5128 4326
rect 5152 4324 5208 4326
rect 5232 4324 5288 4326
rect 5312 4324 5368 4326
rect 5078 4120 5134 4176
rect 7572 11450 7628 11452
rect 7652 11450 7708 11452
rect 7732 11450 7788 11452
rect 7812 11450 7868 11452
rect 7572 11398 7618 11450
rect 7618 11398 7628 11450
rect 7652 11398 7682 11450
rect 7682 11398 7694 11450
rect 7694 11398 7708 11450
rect 7732 11398 7746 11450
rect 7746 11398 7758 11450
rect 7758 11398 7788 11450
rect 7812 11398 7822 11450
rect 7822 11398 7868 11450
rect 7572 11396 7628 11398
rect 7652 11396 7708 11398
rect 7732 11396 7788 11398
rect 7812 11396 7868 11398
rect 5538 5072 5594 5128
rect 5072 3290 5128 3292
rect 5152 3290 5208 3292
rect 5232 3290 5288 3292
rect 5312 3290 5368 3292
rect 5072 3238 5118 3290
rect 5118 3238 5128 3290
rect 5152 3238 5182 3290
rect 5182 3238 5194 3290
rect 5194 3238 5208 3290
rect 5232 3238 5246 3290
rect 5246 3238 5258 3290
rect 5258 3238 5288 3290
rect 5312 3238 5322 3290
rect 5322 3238 5368 3290
rect 5072 3236 5128 3238
rect 5152 3236 5208 3238
rect 5232 3236 5288 3238
rect 5312 3236 5368 3238
rect 6734 10104 6790 10160
rect 6734 9288 6790 9344
rect 6918 6568 6974 6624
rect 6826 5344 6882 5400
rect 7572 10362 7628 10364
rect 7652 10362 7708 10364
rect 7732 10362 7788 10364
rect 7812 10362 7868 10364
rect 7572 10310 7618 10362
rect 7618 10310 7628 10362
rect 7652 10310 7682 10362
rect 7682 10310 7694 10362
rect 7694 10310 7708 10362
rect 7732 10310 7746 10362
rect 7746 10310 7758 10362
rect 7758 10310 7788 10362
rect 7812 10310 7822 10362
rect 7822 10310 7868 10362
rect 7572 10308 7628 10310
rect 7652 10308 7708 10310
rect 7732 10308 7788 10310
rect 7812 10308 7868 10310
rect 8022 10648 8078 10704
rect 7572 9274 7628 9276
rect 7652 9274 7708 9276
rect 7732 9274 7788 9276
rect 7812 9274 7868 9276
rect 7572 9222 7618 9274
rect 7618 9222 7628 9274
rect 7652 9222 7682 9274
rect 7682 9222 7694 9274
rect 7694 9222 7708 9274
rect 7732 9222 7746 9274
rect 7746 9222 7758 9274
rect 7758 9222 7788 9274
rect 7812 9222 7822 9274
rect 7822 9222 7868 9274
rect 7572 9220 7628 9222
rect 7652 9220 7708 9222
rect 7732 9220 7788 9222
rect 7812 9220 7868 9222
rect 7378 9016 7434 9072
rect 7572 8186 7628 8188
rect 7652 8186 7708 8188
rect 7732 8186 7788 8188
rect 7812 8186 7868 8188
rect 7572 8134 7618 8186
rect 7618 8134 7628 8186
rect 7652 8134 7682 8186
rect 7682 8134 7694 8186
rect 7694 8134 7708 8186
rect 7732 8134 7746 8186
rect 7746 8134 7758 8186
rect 7758 8134 7788 8186
rect 7812 8134 7822 8186
rect 7822 8134 7868 8186
rect 7572 8132 7628 8134
rect 7652 8132 7708 8134
rect 7732 8132 7788 8134
rect 7812 8132 7868 8134
rect 7572 7098 7628 7100
rect 7652 7098 7708 7100
rect 7732 7098 7788 7100
rect 7812 7098 7868 7100
rect 7572 7046 7618 7098
rect 7618 7046 7628 7098
rect 7652 7046 7682 7098
rect 7682 7046 7694 7098
rect 7694 7046 7708 7098
rect 7732 7046 7746 7098
rect 7746 7046 7758 7098
rect 7758 7046 7788 7098
rect 7812 7046 7822 7098
rect 7822 7046 7868 7098
rect 7572 7044 7628 7046
rect 7652 7044 7708 7046
rect 7732 7044 7788 7046
rect 7812 7044 7868 7046
rect 8114 6976 8170 7032
rect 7572 6010 7628 6012
rect 7652 6010 7708 6012
rect 7732 6010 7788 6012
rect 7812 6010 7868 6012
rect 7572 5958 7618 6010
rect 7618 5958 7628 6010
rect 7652 5958 7682 6010
rect 7682 5958 7694 6010
rect 7694 5958 7708 6010
rect 7732 5958 7746 6010
rect 7746 5958 7758 6010
rect 7758 5958 7788 6010
rect 7812 5958 7822 6010
rect 7822 5958 7868 6010
rect 7572 5956 7628 5958
rect 7652 5956 7708 5958
rect 7732 5956 7788 5958
rect 7812 5956 7868 5958
rect 7572 4922 7628 4924
rect 7652 4922 7708 4924
rect 7732 4922 7788 4924
rect 7812 4922 7868 4924
rect 7572 4870 7618 4922
rect 7618 4870 7628 4922
rect 7652 4870 7682 4922
rect 7682 4870 7694 4922
rect 7694 4870 7708 4922
rect 7732 4870 7746 4922
rect 7746 4870 7758 4922
rect 7758 4870 7788 4922
rect 7812 4870 7822 4922
rect 7822 4870 7868 4922
rect 7572 4868 7628 4870
rect 7652 4868 7708 4870
rect 7732 4868 7788 4870
rect 7812 4868 7868 4870
rect 7572 3834 7628 3836
rect 7652 3834 7708 3836
rect 7732 3834 7788 3836
rect 7812 3834 7868 3836
rect 7572 3782 7618 3834
rect 7618 3782 7628 3834
rect 7652 3782 7682 3834
rect 7682 3782 7694 3834
rect 7694 3782 7708 3834
rect 7732 3782 7746 3834
rect 7746 3782 7758 3834
rect 7758 3782 7788 3834
rect 7812 3782 7822 3834
rect 7822 3782 7868 3834
rect 7572 3780 7628 3782
rect 7652 3780 7708 3782
rect 7732 3780 7788 3782
rect 7812 3780 7868 3782
rect 7286 3440 7342 3496
rect 6826 3304 6882 3360
rect 5072 2202 5128 2204
rect 5152 2202 5208 2204
rect 5232 2202 5288 2204
rect 5312 2202 5368 2204
rect 5072 2150 5118 2202
rect 5118 2150 5128 2202
rect 5152 2150 5182 2202
rect 5182 2150 5194 2202
rect 5194 2150 5208 2202
rect 5232 2150 5246 2202
rect 5246 2150 5258 2202
rect 5258 2150 5288 2202
rect 5312 2150 5322 2202
rect 5322 2150 5368 2202
rect 5072 2148 5128 2150
rect 5152 2148 5208 2150
rect 5232 2148 5288 2150
rect 5312 2148 5368 2150
rect 6550 2488 6606 2544
rect 9126 8200 9182 8256
rect 16578 11872 16634 11928
rect 20718 11464 20774 11520
rect 16578 11056 16634 11112
rect 16578 9424 16634 9480
rect 16578 8628 16634 8664
rect 16578 8608 16580 8628
rect 16580 8608 16632 8628
rect 16632 8608 16634 8628
rect 9218 7792 9274 7848
rect 16670 7384 16726 7440
rect 9218 6160 9274 6216
rect 8758 4528 8814 4584
rect 8390 2896 8446 2952
rect 7572 2746 7628 2748
rect 7652 2746 7708 2748
rect 7732 2746 7788 2748
rect 7812 2746 7868 2748
rect 7572 2694 7618 2746
rect 7618 2694 7628 2746
rect 7652 2694 7682 2746
rect 7682 2694 7694 2746
rect 7694 2694 7708 2746
rect 7732 2694 7746 2746
rect 7746 2694 7758 2746
rect 7758 2694 7788 2746
rect 7812 2694 7822 2746
rect 7822 2694 7868 2746
rect 7572 2692 7628 2694
rect 7652 2692 7708 2694
rect 7732 2692 7788 2694
rect 7812 2692 7868 2694
rect 9586 5752 9642 5808
rect 7572 1658 7628 1660
rect 7652 1658 7708 1660
rect 7732 1658 7788 1660
rect 7812 1658 7868 1660
rect 7572 1606 7618 1658
rect 7618 1606 7628 1658
rect 7652 1606 7682 1658
rect 7682 1606 7694 1658
rect 7694 1606 7708 1658
rect 7732 1606 7746 1658
rect 7746 1606 7758 1658
rect 7758 1606 7788 1658
rect 7812 1606 7822 1658
rect 7822 1606 7868 1658
rect 7572 1604 7628 1606
rect 7652 1604 7708 1606
rect 7732 1604 7788 1606
rect 7812 1604 7868 1606
rect 5072 1114 5128 1116
rect 5152 1114 5208 1116
rect 5232 1114 5288 1116
rect 5312 1114 5368 1116
rect 5072 1062 5118 1114
rect 5118 1062 5128 1114
rect 5152 1062 5182 1114
rect 5182 1062 5194 1114
rect 5194 1062 5208 1114
rect 5232 1062 5246 1114
rect 5246 1062 5258 1114
rect 5258 1062 5288 1114
rect 5312 1062 5322 1114
rect 5322 1062 5368 1114
rect 5072 1060 5128 1062
rect 5152 1060 5208 1062
rect 5232 1060 5288 1062
rect 5312 1060 5368 1062
rect 9126 856 9182 912
rect 16578 4120 16634 4176
rect 11518 3712 11574 3768
rect 16578 2080 16634 2136
rect 9494 1672 9550 1728
rect 9402 1264 9458 1320
rect 9218 448 9274 504
<< metal3 >>
rect 9489 12338 9555 12341
rect 14000 12338 34000 12368
rect 9489 12336 34000 12338
rect 9489 12280 9494 12336
rect 9550 12280 34000 12336
rect 9489 12278 34000 12280
rect 9489 12275 9555 12278
rect 14000 12248 34000 12278
rect 14000 11928 34000 11960
rect 14000 11872 16578 11928
rect 16634 11872 34000 11928
rect 14000 11840 34000 11872
rect 14000 11520 34000 11552
rect 14000 11464 20718 11520
rect 20774 11464 34000 11520
rect 2560 11456 2880 11457
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 11391 2880 11392
rect 7560 11456 7880 11457
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 14000 11432 34000 11464
rect 7560 11391 7880 11392
rect 14000 11112 34000 11144
rect 14000 11056 16578 11112
rect 16634 11056 34000 11112
rect 14000 11024 34000 11056
rect 5060 10912 5380 10913
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 10847 5380 10848
rect 8017 10706 8083 10709
rect 14000 10706 34000 10736
rect 8017 10704 34000 10706
rect 8017 10648 8022 10704
rect 8078 10648 34000 10704
rect 8017 10646 34000 10648
rect 8017 10643 8083 10646
rect 14000 10616 34000 10646
rect 2560 10368 2880 10369
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 10303 2880 10304
rect 7560 10368 7880 10369
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 10303 7880 10304
rect 14000 10298 34000 10328
rect 12390 10238 34000 10298
rect 6729 10162 6795 10165
rect 12390 10162 12450 10238
rect 14000 10208 34000 10238
rect 6729 10160 12450 10162
rect 6729 10104 6734 10160
rect 6790 10104 12450 10160
rect 6729 10102 12450 10104
rect 6729 10099 6795 10102
rect 1485 10026 1551 10029
rect 1485 10024 12450 10026
rect 1485 9968 1490 10024
rect 1546 9968 12450 10024
rect 1485 9966 12450 9968
rect 1485 9963 1551 9966
rect 12390 9890 12450 9966
rect 14000 9890 34000 9920
rect 12390 9830 34000 9890
rect 5060 9824 5380 9825
rect 5060 9760 5068 9824
rect 5132 9760 5148 9824
rect 5212 9760 5228 9824
rect 5292 9760 5308 9824
rect 5372 9760 5380 9824
rect 14000 9800 34000 9830
rect 5060 9759 5380 9760
rect 3233 9482 3299 9485
rect 4705 9482 4771 9485
rect 3233 9480 4771 9482
rect 3233 9424 3238 9480
rect 3294 9424 4710 9480
rect 4766 9424 4771 9480
rect 3233 9422 4771 9424
rect 3233 9419 3299 9422
rect 4705 9419 4771 9422
rect 14000 9480 34000 9512
rect 14000 9424 16578 9480
rect 16634 9424 34000 9480
rect 14000 9392 34000 9424
rect 5993 9346 6059 9349
rect 6729 9346 6795 9349
rect 5993 9344 6795 9346
rect 5993 9288 5998 9344
rect 6054 9288 6734 9344
rect 6790 9288 6795 9344
rect 5993 9286 6795 9288
rect 5993 9283 6059 9286
rect 6729 9283 6795 9286
rect 2560 9280 2880 9281
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 9215 2880 9216
rect 7560 9280 7880 9281
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 9215 7880 9216
rect 7373 9074 7439 9077
rect 14000 9074 34000 9104
rect 7373 9072 34000 9074
rect 7373 9016 7378 9072
rect 7434 9016 34000 9072
rect 7373 9014 34000 9016
rect 7373 9011 7439 9014
rect 14000 8984 34000 9014
rect 5060 8736 5380 8737
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 8671 5380 8672
rect 14000 8664 34000 8696
rect 14000 8608 16578 8664
rect 16634 8608 34000 8664
rect 14000 8576 34000 8608
rect 9121 8258 9187 8261
rect 14000 8258 34000 8288
rect 9121 8256 34000 8258
rect 9121 8200 9126 8256
rect 9182 8200 34000 8256
rect 9121 8198 34000 8200
rect 9121 8195 9187 8198
rect 2560 8192 2880 8193
rect 2560 8128 2568 8192
rect 2632 8128 2648 8192
rect 2712 8128 2728 8192
rect 2792 8128 2808 8192
rect 2872 8128 2880 8192
rect 2560 8127 2880 8128
rect 7560 8192 7880 8193
rect 7560 8128 7568 8192
rect 7632 8128 7648 8192
rect 7712 8128 7728 8192
rect 7792 8128 7808 8192
rect 7872 8128 7880 8192
rect 14000 8168 34000 8198
rect 7560 8127 7880 8128
rect 9213 7850 9279 7853
rect 14000 7850 34000 7880
rect 9213 7848 34000 7850
rect 9213 7792 9218 7848
rect 9274 7792 34000 7848
rect 9213 7790 34000 7792
rect 9213 7787 9279 7790
rect 14000 7760 34000 7790
rect 5060 7648 5380 7649
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 7583 5380 7584
rect 14000 7440 34000 7472
rect 14000 7384 16670 7440
rect 16726 7384 34000 7440
rect 14000 7352 34000 7384
rect 2560 7104 2880 7105
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 7039 2880 7040
rect 7560 7104 7880 7105
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 7039 7880 7040
rect 8109 7034 8175 7037
rect 14000 7034 34000 7064
rect 8109 7032 34000 7034
rect 8109 6976 8114 7032
rect 8170 6976 34000 7032
rect 8109 6974 34000 6976
rect 8109 6971 8175 6974
rect 14000 6944 34000 6974
rect 6913 6626 6979 6629
rect 14000 6626 34000 6656
rect 6913 6624 34000 6626
rect 6913 6568 6918 6624
rect 6974 6568 34000 6624
rect 6913 6566 34000 6568
rect 6913 6563 6979 6566
rect 5060 6560 5380 6561
rect 5060 6496 5068 6560
rect 5132 6496 5148 6560
rect 5212 6496 5228 6560
rect 5292 6496 5308 6560
rect 5372 6496 5380 6560
rect 14000 6536 34000 6566
rect 5060 6495 5380 6496
rect 9213 6218 9279 6221
rect 14000 6218 34000 6248
rect 9213 6216 34000 6218
rect 9213 6160 9218 6216
rect 9274 6160 34000 6216
rect 9213 6158 34000 6160
rect 9213 6155 9279 6158
rect 14000 6128 34000 6158
rect 2560 6016 2880 6017
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 5951 2880 5952
rect 7560 6016 7880 6017
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 5951 7880 5952
rect 9581 5810 9647 5813
rect 14000 5810 34000 5840
rect 9581 5808 34000 5810
rect 9581 5752 9586 5808
rect 9642 5752 34000 5808
rect 9581 5750 34000 5752
rect 9581 5747 9647 5750
rect 14000 5720 34000 5750
rect 5060 5472 5380 5473
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 5407 5380 5408
rect 6821 5402 6887 5405
rect 14000 5402 34000 5432
rect 6821 5400 34000 5402
rect 6821 5344 6826 5400
rect 6882 5344 34000 5400
rect 6821 5342 34000 5344
rect 6821 5339 6887 5342
rect 14000 5312 34000 5342
rect 5533 5130 5599 5133
rect 5533 5128 12450 5130
rect 5533 5072 5538 5128
rect 5594 5072 12450 5128
rect 5533 5070 12450 5072
rect 5533 5067 5599 5070
rect 12390 4994 12450 5070
rect 14000 4994 34000 5024
rect 12390 4934 34000 4994
rect 7560 4928 7880 4929
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 14000 4904 34000 4934
rect 7560 4863 7880 4864
rect 8753 4586 8819 4589
rect 14000 4586 34000 4616
rect 8753 4584 34000 4586
rect 8753 4528 8758 4584
rect 8814 4528 34000 4584
rect 8753 4526 34000 4528
rect 8753 4523 8819 4526
rect 14000 4496 34000 4526
rect 5060 4384 5380 4385
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 4319 5380 4320
rect 4705 4312 4771 4317
rect 4705 4256 4710 4312
rect 4766 4256 4771 4312
rect 4705 4251 4771 4256
rect 4708 4178 4768 4251
rect 5073 4178 5139 4181
rect 4708 4176 5139 4178
rect 4708 4120 5078 4176
rect 5134 4120 5139 4176
rect 4708 4118 5139 4120
rect 5073 4115 5139 4118
rect 14000 4176 34000 4208
rect 14000 4120 16578 4176
rect 16634 4120 34000 4176
rect 14000 4088 34000 4120
rect 7560 3840 7880 3841
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 3775 7880 3776
rect 11513 3770 11579 3773
rect 14000 3770 34000 3800
rect 11513 3768 34000 3770
rect 11513 3712 11518 3768
rect 11574 3712 34000 3768
rect 11513 3710 34000 3712
rect 11513 3707 11579 3710
rect 14000 3680 34000 3710
rect 3417 3498 3483 3501
rect 7281 3498 7347 3501
rect 3417 3496 7347 3498
rect 3417 3440 3422 3496
rect 3478 3440 7286 3496
rect 7342 3440 7347 3496
rect 3417 3438 7347 3440
rect 3417 3435 3483 3438
rect 7281 3435 7347 3438
rect 2681 3362 2747 3365
rect 2484 3360 2747 3362
rect 2484 3304 2686 3360
rect 2742 3304 2747 3360
rect 2484 3302 2747 3304
rect 2681 3299 2747 3302
rect 6821 3362 6887 3365
rect 14000 3362 34000 3392
rect 6821 3360 34000 3362
rect 6821 3304 6826 3360
rect 6882 3304 34000 3360
rect 6821 3302 34000 3304
rect 6821 3299 6887 3302
rect 5060 3296 5380 3297
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 14000 3272 34000 3302
rect 5060 3231 5380 3232
rect 8385 2954 8451 2957
rect 14000 2954 34000 2984
rect 8385 2952 34000 2954
rect 8385 2896 8390 2952
rect 8446 2896 34000 2952
rect 8385 2894 34000 2896
rect 8385 2891 8451 2894
rect 14000 2864 34000 2894
rect 7560 2752 7880 2753
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 2687 7880 2688
rect 6545 2546 6611 2549
rect 14000 2546 34000 2576
rect 6545 2544 34000 2546
rect 6545 2488 6550 2544
rect 6606 2488 34000 2544
rect 6545 2486 34000 2488
rect 6545 2483 6611 2486
rect 14000 2456 34000 2486
rect 5060 2208 5380 2209
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 2143 5380 2144
rect 14000 2136 34000 2168
rect 14000 2080 16578 2136
rect 16634 2080 34000 2136
rect 14000 2048 34000 2080
rect 9489 1730 9555 1733
rect 14000 1730 34000 1760
rect 9489 1728 34000 1730
rect 9489 1672 9494 1728
rect 9550 1672 34000 1728
rect 9489 1670 34000 1672
rect 9489 1667 9555 1670
rect 7560 1664 7880 1665
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 14000 1640 34000 1670
rect 7560 1599 7880 1600
rect 9397 1322 9463 1325
rect 14000 1322 34000 1352
rect 9397 1320 34000 1322
rect 9397 1264 9402 1320
rect 9458 1264 34000 1320
rect 9397 1262 34000 1264
rect 9397 1259 9463 1262
rect 14000 1232 34000 1262
rect 5060 1120 5380 1121
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 5060 1055 5380 1056
rect 9121 914 9187 917
rect 14000 914 34000 944
rect 9121 912 34000 914
rect 9121 856 9126 912
rect 9182 856 34000 912
rect 9121 854 34000 856
rect 9121 851 9187 854
rect 14000 824 34000 854
rect 9213 506 9279 509
rect 14000 506 34000 536
rect 9213 504 34000 506
rect 9213 448 9218 504
rect 9274 448 34000 504
rect 9213 446 34000 448
rect 9213 443 9279 446
rect 14000 416 34000 446
<< via3 >>
rect 2568 11452 2632 11456
rect 2568 11396 2572 11452
rect 2572 11396 2628 11452
rect 2628 11396 2632 11452
rect 2568 11392 2632 11396
rect 2648 11452 2712 11456
rect 2648 11396 2652 11452
rect 2652 11396 2708 11452
rect 2708 11396 2712 11452
rect 2648 11392 2712 11396
rect 2728 11452 2792 11456
rect 2728 11396 2732 11452
rect 2732 11396 2788 11452
rect 2788 11396 2792 11452
rect 2728 11392 2792 11396
rect 2808 11452 2872 11456
rect 2808 11396 2812 11452
rect 2812 11396 2868 11452
rect 2868 11396 2872 11452
rect 2808 11392 2872 11396
rect 7568 11452 7632 11456
rect 7568 11396 7572 11452
rect 7572 11396 7628 11452
rect 7628 11396 7632 11452
rect 7568 11392 7632 11396
rect 7648 11452 7712 11456
rect 7648 11396 7652 11452
rect 7652 11396 7708 11452
rect 7708 11396 7712 11452
rect 7648 11392 7712 11396
rect 7728 11452 7792 11456
rect 7728 11396 7732 11452
rect 7732 11396 7788 11452
rect 7788 11396 7792 11452
rect 7728 11392 7792 11396
rect 7808 11452 7872 11456
rect 7808 11396 7812 11452
rect 7812 11396 7868 11452
rect 7868 11396 7872 11452
rect 7808 11392 7872 11396
rect 5068 10908 5132 10912
rect 5068 10852 5072 10908
rect 5072 10852 5128 10908
rect 5128 10852 5132 10908
rect 5068 10848 5132 10852
rect 5148 10908 5212 10912
rect 5148 10852 5152 10908
rect 5152 10852 5208 10908
rect 5208 10852 5212 10908
rect 5148 10848 5212 10852
rect 5228 10908 5292 10912
rect 5228 10852 5232 10908
rect 5232 10852 5288 10908
rect 5288 10852 5292 10908
rect 5228 10848 5292 10852
rect 5308 10908 5372 10912
rect 5308 10852 5312 10908
rect 5312 10852 5368 10908
rect 5368 10852 5372 10908
rect 5308 10848 5372 10852
rect 2568 10364 2632 10368
rect 2568 10308 2572 10364
rect 2572 10308 2628 10364
rect 2628 10308 2632 10364
rect 2568 10304 2632 10308
rect 2648 10364 2712 10368
rect 2648 10308 2652 10364
rect 2652 10308 2708 10364
rect 2708 10308 2712 10364
rect 2648 10304 2712 10308
rect 2728 10364 2792 10368
rect 2728 10308 2732 10364
rect 2732 10308 2788 10364
rect 2788 10308 2792 10364
rect 2728 10304 2792 10308
rect 2808 10364 2872 10368
rect 2808 10308 2812 10364
rect 2812 10308 2868 10364
rect 2868 10308 2872 10364
rect 2808 10304 2872 10308
rect 7568 10364 7632 10368
rect 7568 10308 7572 10364
rect 7572 10308 7628 10364
rect 7628 10308 7632 10364
rect 7568 10304 7632 10308
rect 7648 10364 7712 10368
rect 7648 10308 7652 10364
rect 7652 10308 7708 10364
rect 7708 10308 7712 10364
rect 7648 10304 7712 10308
rect 7728 10364 7792 10368
rect 7728 10308 7732 10364
rect 7732 10308 7788 10364
rect 7788 10308 7792 10364
rect 7728 10304 7792 10308
rect 7808 10364 7872 10368
rect 7808 10308 7812 10364
rect 7812 10308 7868 10364
rect 7868 10308 7872 10364
rect 7808 10304 7872 10308
rect 5068 9820 5132 9824
rect 5068 9764 5072 9820
rect 5072 9764 5128 9820
rect 5128 9764 5132 9820
rect 5068 9760 5132 9764
rect 5148 9820 5212 9824
rect 5148 9764 5152 9820
rect 5152 9764 5208 9820
rect 5208 9764 5212 9820
rect 5148 9760 5212 9764
rect 5228 9820 5292 9824
rect 5228 9764 5232 9820
rect 5232 9764 5288 9820
rect 5288 9764 5292 9820
rect 5228 9760 5292 9764
rect 5308 9820 5372 9824
rect 5308 9764 5312 9820
rect 5312 9764 5368 9820
rect 5368 9764 5372 9820
rect 5308 9760 5372 9764
rect 2568 9276 2632 9280
rect 2568 9220 2572 9276
rect 2572 9220 2628 9276
rect 2628 9220 2632 9276
rect 2568 9216 2632 9220
rect 2648 9276 2712 9280
rect 2648 9220 2652 9276
rect 2652 9220 2708 9276
rect 2708 9220 2712 9276
rect 2648 9216 2712 9220
rect 2728 9276 2792 9280
rect 2728 9220 2732 9276
rect 2732 9220 2788 9276
rect 2788 9220 2792 9276
rect 2728 9216 2792 9220
rect 2808 9276 2872 9280
rect 2808 9220 2812 9276
rect 2812 9220 2868 9276
rect 2868 9220 2872 9276
rect 2808 9216 2872 9220
rect 7568 9276 7632 9280
rect 7568 9220 7572 9276
rect 7572 9220 7628 9276
rect 7628 9220 7632 9276
rect 7568 9216 7632 9220
rect 7648 9276 7712 9280
rect 7648 9220 7652 9276
rect 7652 9220 7708 9276
rect 7708 9220 7712 9276
rect 7648 9216 7712 9220
rect 7728 9276 7792 9280
rect 7728 9220 7732 9276
rect 7732 9220 7788 9276
rect 7788 9220 7792 9276
rect 7728 9216 7792 9220
rect 7808 9276 7872 9280
rect 7808 9220 7812 9276
rect 7812 9220 7868 9276
rect 7868 9220 7872 9276
rect 7808 9216 7872 9220
rect 5068 8732 5132 8736
rect 5068 8676 5072 8732
rect 5072 8676 5128 8732
rect 5128 8676 5132 8732
rect 5068 8672 5132 8676
rect 5148 8732 5212 8736
rect 5148 8676 5152 8732
rect 5152 8676 5208 8732
rect 5208 8676 5212 8732
rect 5148 8672 5212 8676
rect 5228 8732 5292 8736
rect 5228 8676 5232 8732
rect 5232 8676 5288 8732
rect 5288 8676 5292 8732
rect 5228 8672 5292 8676
rect 5308 8732 5372 8736
rect 5308 8676 5312 8732
rect 5312 8676 5368 8732
rect 5368 8676 5372 8732
rect 5308 8672 5372 8676
rect 2568 8188 2632 8192
rect 2568 8132 2572 8188
rect 2572 8132 2628 8188
rect 2628 8132 2632 8188
rect 2568 8128 2632 8132
rect 2648 8188 2712 8192
rect 2648 8132 2652 8188
rect 2652 8132 2708 8188
rect 2708 8132 2712 8188
rect 2648 8128 2712 8132
rect 2728 8188 2792 8192
rect 2728 8132 2732 8188
rect 2732 8132 2788 8188
rect 2788 8132 2792 8188
rect 2728 8128 2792 8132
rect 2808 8188 2872 8192
rect 2808 8132 2812 8188
rect 2812 8132 2868 8188
rect 2868 8132 2872 8188
rect 2808 8128 2872 8132
rect 7568 8188 7632 8192
rect 7568 8132 7572 8188
rect 7572 8132 7628 8188
rect 7628 8132 7632 8188
rect 7568 8128 7632 8132
rect 7648 8188 7712 8192
rect 7648 8132 7652 8188
rect 7652 8132 7708 8188
rect 7708 8132 7712 8188
rect 7648 8128 7712 8132
rect 7728 8188 7792 8192
rect 7728 8132 7732 8188
rect 7732 8132 7788 8188
rect 7788 8132 7792 8188
rect 7728 8128 7792 8132
rect 7808 8188 7872 8192
rect 7808 8132 7812 8188
rect 7812 8132 7868 8188
rect 7868 8132 7872 8188
rect 7808 8128 7872 8132
rect 5068 7644 5132 7648
rect 5068 7588 5072 7644
rect 5072 7588 5128 7644
rect 5128 7588 5132 7644
rect 5068 7584 5132 7588
rect 5148 7644 5212 7648
rect 5148 7588 5152 7644
rect 5152 7588 5208 7644
rect 5208 7588 5212 7644
rect 5148 7584 5212 7588
rect 5228 7644 5292 7648
rect 5228 7588 5232 7644
rect 5232 7588 5288 7644
rect 5288 7588 5292 7644
rect 5228 7584 5292 7588
rect 5308 7644 5372 7648
rect 5308 7588 5312 7644
rect 5312 7588 5368 7644
rect 5368 7588 5372 7644
rect 5308 7584 5372 7588
rect 2568 7100 2632 7104
rect 2568 7044 2572 7100
rect 2572 7044 2628 7100
rect 2628 7044 2632 7100
rect 2568 7040 2632 7044
rect 2648 7100 2712 7104
rect 2648 7044 2652 7100
rect 2652 7044 2708 7100
rect 2708 7044 2712 7100
rect 2648 7040 2712 7044
rect 2728 7100 2792 7104
rect 2728 7044 2732 7100
rect 2732 7044 2788 7100
rect 2788 7044 2792 7100
rect 2728 7040 2792 7044
rect 2808 7100 2872 7104
rect 2808 7044 2812 7100
rect 2812 7044 2868 7100
rect 2868 7044 2872 7100
rect 2808 7040 2872 7044
rect 7568 7100 7632 7104
rect 7568 7044 7572 7100
rect 7572 7044 7628 7100
rect 7628 7044 7632 7100
rect 7568 7040 7632 7044
rect 7648 7100 7712 7104
rect 7648 7044 7652 7100
rect 7652 7044 7708 7100
rect 7708 7044 7712 7100
rect 7648 7040 7712 7044
rect 7728 7100 7792 7104
rect 7728 7044 7732 7100
rect 7732 7044 7788 7100
rect 7788 7044 7792 7100
rect 7728 7040 7792 7044
rect 7808 7100 7872 7104
rect 7808 7044 7812 7100
rect 7812 7044 7868 7100
rect 7868 7044 7872 7100
rect 7808 7040 7872 7044
rect 5068 6556 5132 6560
rect 5068 6500 5072 6556
rect 5072 6500 5128 6556
rect 5128 6500 5132 6556
rect 5068 6496 5132 6500
rect 5148 6556 5212 6560
rect 5148 6500 5152 6556
rect 5152 6500 5208 6556
rect 5208 6500 5212 6556
rect 5148 6496 5212 6500
rect 5228 6556 5292 6560
rect 5228 6500 5232 6556
rect 5232 6500 5288 6556
rect 5288 6500 5292 6556
rect 5228 6496 5292 6500
rect 5308 6556 5372 6560
rect 5308 6500 5312 6556
rect 5312 6500 5368 6556
rect 5368 6500 5372 6556
rect 5308 6496 5372 6500
rect 2568 6012 2632 6016
rect 2568 5956 2572 6012
rect 2572 5956 2628 6012
rect 2628 5956 2632 6012
rect 2568 5952 2632 5956
rect 2648 6012 2712 6016
rect 2648 5956 2652 6012
rect 2652 5956 2708 6012
rect 2708 5956 2712 6012
rect 2648 5952 2712 5956
rect 2728 6012 2792 6016
rect 2728 5956 2732 6012
rect 2732 5956 2788 6012
rect 2788 5956 2792 6012
rect 2728 5952 2792 5956
rect 2808 6012 2872 6016
rect 2808 5956 2812 6012
rect 2812 5956 2868 6012
rect 2868 5956 2872 6012
rect 2808 5952 2872 5956
rect 7568 6012 7632 6016
rect 7568 5956 7572 6012
rect 7572 5956 7628 6012
rect 7628 5956 7632 6012
rect 7568 5952 7632 5956
rect 7648 6012 7712 6016
rect 7648 5956 7652 6012
rect 7652 5956 7708 6012
rect 7708 5956 7712 6012
rect 7648 5952 7712 5956
rect 7728 6012 7792 6016
rect 7728 5956 7732 6012
rect 7732 5956 7788 6012
rect 7788 5956 7792 6012
rect 7728 5952 7792 5956
rect 7808 6012 7872 6016
rect 7808 5956 7812 6012
rect 7812 5956 7868 6012
rect 7868 5956 7872 6012
rect 7808 5952 7872 5956
rect 5068 5468 5132 5472
rect 5068 5412 5072 5468
rect 5072 5412 5128 5468
rect 5128 5412 5132 5468
rect 5068 5408 5132 5412
rect 5148 5468 5212 5472
rect 5148 5412 5152 5468
rect 5152 5412 5208 5468
rect 5208 5412 5212 5468
rect 5148 5408 5212 5412
rect 5228 5468 5292 5472
rect 5228 5412 5232 5468
rect 5232 5412 5288 5468
rect 5288 5412 5292 5468
rect 5228 5408 5292 5412
rect 5308 5468 5372 5472
rect 5308 5412 5312 5468
rect 5312 5412 5368 5468
rect 5368 5412 5372 5468
rect 5308 5408 5372 5412
rect 7568 4924 7632 4928
rect 7568 4868 7572 4924
rect 7572 4868 7628 4924
rect 7628 4868 7632 4924
rect 7568 4864 7632 4868
rect 7648 4924 7712 4928
rect 7648 4868 7652 4924
rect 7652 4868 7708 4924
rect 7708 4868 7712 4924
rect 7648 4864 7712 4868
rect 7728 4924 7792 4928
rect 7728 4868 7732 4924
rect 7732 4868 7788 4924
rect 7788 4868 7792 4924
rect 7728 4864 7792 4868
rect 7808 4924 7872 4928
rect 7808 4868 7812 4924
rect 7812 4868 7868 4924
rect 7868 4868 7872 4924
rect 7808 4864 7872 4868
rect 5068 4380 5132 4384
rect 5068 4324 5072 4380
rect 5072 4324 5128 4380
rect 5128 4324 5132 4380
rect 5068 4320 5132 4324
rect 5148 4380 5212 4384
rect 5148 4324 5152 4380
rect 5152 4324 5208 4380
rect 5208 4324 5212 4380
rect 5148 4320 5212 4324
rect 5228 4380 5292 4384
rect 5228 4324 5232 4380
rect 5232 4324 5288 4380
rect 5288 4324 5292 4380
rect 5228 4320 5292 4324
rect 5308 4380 5372 4384
rect 5308 4324 5312 4380
rect 5312 4324 5368 4380
rect 5368 4324 5372 4380
rect 5308 4320 5372 4324
rect 7568 3836 7632 3840
rect 7568 3780 7572 3836
rect 7572 3780 7628 3836
rect 7628 3780 7632 3836
rect 7568 3776 7632 3780
rect 7648 3836 7712 3840
rect 7648 3780 7652 3836
rect 7652 3780 7708 3836
rect 7708 3780 7712 3836
rect 7648 3776 7712 3780
rect 7728 3836 7792 3840
rect 7728 3780 7732 3836
rect 7732 3780 7788 3836
rect 7788 3780 7792 3836
rect 7728 3776 7792 3780
rect 7808 3836 7872 3840
rect 7808 3780 7812 3836
rect 7812 3780 7868 3836
rect 7868 3780 7872 3836
rect 7808 3776 7872 3780
rect 5068 3292 5132 3296
rect 5068 3236 5072 3292
rect 5072 3236 5128 3292
rect 5128 3236 5132 3292
rect 5068 3232 5132 3236
rect 5148 3292 5212 3296
rect 5148 3236 5152 3292
rect 5152 3236 5208 3292
rect 5208 3236 5212 3292
rect 5148 3232 5212 3236
rect 5228 3292 5292 3296
rect 5228 3236 5232 3292
rect 5232 3236 5288 3292
rect 5288 3236 5292 3292
rect 5228 3232 5292 3236
rect 5308 3292 5372 3296
rect 5308 3236 5312 3292
rect 5312 3236 5368 3292
rect 5368 3236 5372 3292
rect 5308 3232 5372 3236
rect 7568 2748 7632 2752
rect 7568 2692 7572 2748
rect 7572 2692 7628 2748
rect 7628 2692 7632 2748
rect 7568 2688 7632 2692
rect 7648 2748 7712 2752
rect 7648 2692 7652 2748
rect 7652 2692 7708 2748
rect 7708 2692 7712 2748
rect 7648 2688 7712 2692
rect 7728 2748 7792 2752
rect 7728 2692 7732 2748
rect 7732 2692 7788 2748
rect 7788 2692 7792 2748
rect 7728 2688 7792 2692
rect 7808 2748 7872 2752
rect 7808 2692 7812 2748
rect 7812 2692 7868 2748
rect 7868 2692 7872 2748
rect 7808 2688 7872 2692
rect 5068 2204 5132 2208
rect 5068 2148 5072 2204
rect 5072 2148 5128 2204
rect 5128 2148 5132 2204
rect 5068 2144 5132 2148
rect 5148 2204 5212 2208
rect 5148 2148 5152 2204
rect 5152 2148 5208 2204
rect 5208 2148 5212 2204
rect 5148 2144 5212 2148
rect 5228 2204 5292 2208
rect 5228 2148 5232 2204
rect 5232 2148 5288 2204
rect 5288 2148 5292 2204
rect 5228 2144 5292 2148
rect 5308 2204 5372 2208
rect 5308 2148 5312 2204
rect 5312 2148 5368 2204
rect 5368 2148 5372 2204
rect 5308 2144 5372 2148
rect 7568 1660 7632 1664
rect 7568 1604 7572 1660
rect 7572 1604 7628 1660
rect 7628 1604 7632 1660
rect 7568 1600 7632 1604
rect 7648 1660 7712 1664
rect 7648 1604 7652 1660
rect 7652 1604 7708 1660
rect 7708 1604 7712 1660
rect 7648 1600 7712 1604
rect 7728 1660 7792 1664
rect 7728 1604 7732 1660
rect 7732 1604 7788 1660
rect 7788 1604 7792 1660
rect 7728 1600 7792 1604
rect 7808 1660 7872 1664
rect 7808 1604 7812 1660
rect 7812 1604 7868 1660
rect 7868 1604 7872 1660
rect 7808 1600 7872 1604
rect 5068 1116 5132 1120
rect 5068 1060 5072 1116
rect 5072 1060 5128 1116
rect 5128 1060 5132 1116
rect 5068 1056 5132 1060
rect 5148 1116 5212 1120
rect 5148 1060 5152 1116
rect 5152 1060 5208 1116
rect 5208 1060 5212 1116
rect 5148 1056 5212 1060
rect 5228 1116 5292 1120
rect 5228 1060 5232 1116
rect 5232 1060 5288 1116
rect 5288 1060 5292 1116
rect 5228 1056 5292 1060
rect 5308 1116 5372 1120
rect 5308 1060 5312 1116
rect 5312 1060 5368 1116
rect 5368 1060 5372 1116
rect 5308 1056 5372 1060
<< metal4 >>
rect 2560 11456 2880 11472
rect 2560 11392 2568 11456
rect 2632 11392 2648 11456
rect 2712 11392 2728 11456
rect 2792 11392 2808 11456
rect 2872 11392 2880 11456
rect 2560 10368 2880 11392
rect 2560 10304 2568 10368
rect 2632 10304 2648 10368
rect 2712 10304 2728 10368
rect 2792 10304 2808 10368
rect 2872 10304 2880 10368
rect 2560 9280 2880 10304
rect 2560 9216 2568 9280
rect 2632 9216 2648 9280
rect 2712 9216 2728 9280
rect 2792 9216 2808 9280
rect 2872 9216 2880 9280
rect 2560 8218 2880 9216
rect 2560 8192 2602 8218
rect 2838 8192 2880 8218
rect 2560 8128 2568 8192
rect 2872 8128 2880 8192
rect 2560 7982 2602 8128
rect 2838 7982 2880 8128
rect 2560 7104 2880 7982
rect 2560 7040 2568 7104
rect 2632 7040 2648 7104
rect 2712 7040 2728 7104
rect 2792 7040 2808 7104
rect 2872 7040 2880 7104
rect 2560 6016 2880 7040
rect 2560 5952 2568 6016
rect 2632 5952 2648 6016
rect 2712 5952 2728 6016
rect 2792 5952 2808 6016
rect 2872 5952 2880 6016
rect 2560 4838 2880 5952
rect 2560 4602 2602 4838
rect 2838 4602 2880 4838
rect 1996 4196 2276 4238
rect 1996 3960 2018 4196
rect 2254 3960 2276 4196
rect 1996 3918 2276 3960
rect 1256 2506 1536 2548
rect 1256 2270 1278 2506
rect 1514 2270 1536 2506
rect 1256 2228 1536 2270
rect 2560 1458 2880 4602
rect 2560 1222 2602 1458
rect 2838 1222 2880 1458
rect 2560 1088 2880 1222
rect 3560 9266 3880 11424
rect 3560 9030 3602 9266
rect 3838 9030 3880 9266
rect 3560 5886 3880 9030
rect 3560 5650 3602 5886
rect 3838 5650 3880 5886
rect 3560 2506 3880 5650
rect 3560 2270 3602 2506
rect 3838 2270 3880 2506
rect 3560 1088 3880 2270
rect 5060 10912 5380 11472
rect 7560 11456 7880 11472
rect 5060 10848 5068 10912
rect 5132 10848 5148 10912
rect 5212 10848 5228 10912
rect 5292 10848 5308 10912
rect 5372 10848 5380 10912
rect 5060 9908 5380 10848
rect 5060 9824 5102 9908
rect 5338 9824 5380 9908
rect 5060 9760 5068 9824
rect 5372 9760 5380 9824
rect 5060 9672 5102 9760
rect 5338 9672 5380 9760
rect 5060 8736 5380 9672
rect 5060 8672 5068 8736
rect 5132 8672 5148 8736
rect 5212 8672 5228 8736
rect 5292 8672 5308 8736
rect 5372 8672 5380 8736
rect 5060 7648 5380 8672
rect 5060 7584 5068 7648
rect 5132 7584 5148 7648
rect 5212 7584 5228 7648
rect 5292 7584 5308 7648
rect 5372 7584 5380 7648
rect 5060 6560 5380 7584
rect 5060 6496 5068 6560
rect 5132 6528 5148 6560
rect 5212 6528 5228 6560
rect 5292 6528 5308 6560
rect 5372 6496 5380 6560
rect 5060 6292 5102 6496
rect 5338 6292 5380 6496
rect 5060 5472 5380 6292
rect 5060 5408 5068 5472
rect 5132 5408 5148 5472
rect 5212 5408 5228 5472
rect 5292 5408 5308 5472
rect 5372 5408 5380 5472
rect 5060 4384 5380 5408
rect 5060 4320 5068 4384
rect 5132 4320 5148 4384
rect 5212 4320 5228 4384
rect 5292 4320 5308 4384
rect 5372 4320 5380 4384
rect 5060 3296 5380 4320
rect 5060 3232 5068 3296
rect 5132 3232 5148 3296
rect 5212 3232 5228 3296
rect 5292 3232 5308 3296
rect 5372 3232 5380 3296
rect 5060 3148 5380 3232
rect 5060 2912 5102 3148
rect 5338 2912 5380 3148
rect 5060 2208 5380 2912
rect 5060 2144 5068 2208
rect 5132 2144 5148 2208
rect 5212 2144 5228 2208
rect 5292 2144 5308 2208
rect 5372 2144 5380 2208
rect 5060 1120 5380 2144
rect 5060 1056 5068 1120
rect 5132 1056 5148 1120
rect 5212 1056 5228 1120
rect 5292 1056 5308 1120
rect 5372 1056 5380 1120
rect 6060 10956 6380 11424
rect 6060 10720 6102 10956
rect 6338 10720 6380 10956
rect 6060 7576 6380 10720
rect 6060 7340 6102 7576
rect 6338 7340 6380 7576
rect 6060 4196 6380 7340
rect 6060 3960 6102 4196
rect 6338 3960 6380 4196
rect 6060 1088 6380 3960
rect 7560 11392 7568 11456
rect 7632 11392 7648 11456
rect 7712 11392 7728 11456
rect 7792 11392 7808 11456
rect 7872 11392 7880 11456
rect 7560 10368 7880 11392
rect 7560 10304 7568 10368
rect 7632 10304 7648 10368
rect 7712 10304 7728 10368
rect 7792 10304 7808 10368
rect 7872 10304 7880 10368
rect 7560 9280 7880 10304
rect 7560 9216 7568 9280
rect 7632 9216 7648 9280
rect 7712 9216 7728 9280
rect 7792 9216 7808 9280
rect 7872 9216 7880 9280
rect 7560 8218 7880 9216
rect 7560 8192 7602 8218
rect 7838 8192 7880 8218
rect 7560 8128 7568 8192
rect 7872 8128 7880 8192
rect 7560 7982 7602 8128
rect 7838 7982 7880 8128
rect 7560 7104 7880 7982
rect 7560 7040 7568 7104
rect 7632 7040 7648 7104
rect 7712 7040 7728 7104
rect 7792 7040 7808 7104
rect 7872 7040 7880 7104
rect 7560 6016 7880 7040
rect 7560 5952 7568 6016
rect 7632 5952 7648 6016
rect 7712 5952 7728 6016
rect 7792 5952 7808 6016
rect 7872 5952 7880 6016
rect 7560 4928 7880 5952
rect 7560 4864 7568 4928
rect 7632 4864 7648 4928
rect 7712 4864 7728 4928
rect 7792 4864 7808 4928
rect 7872 4864 7880 4928
rect 7560 4838 7880 4864
rect 7560 4602 7602 4838
rect 7838 4602 7880 4838
rect 7560 3840 7880 4602
rect 7560 3776 7568 3840
rect 7632 3776 7648 3840
rect 7712 3776 7728 3840
rect 7792 3776 7808 3840
rect 7872 3776 7880 3840
rect 7560 2752 7880 3776
rect 7560 2688 7568 2752
rect 7632 2688 7648 2752
rect 7712 2688 7728 2752
rect 7792 2688 7808 2752
rect 7872 2688 7880 2752
rect 7560 1664 7880 2688
rect 7560 1600 7568 1664
rect 7632 1600 7648 1664
rect 7712 1600 7728 1664
rect 7792 1600 7808 1664
rect 7872 1600 7880 1664
rect 7560 1458 7880 1600
rect 7560 1222 7602 1458
rect 7838 1222 7880 1458
rect 5060 1040 5380 1056
rect 7560 1040 7880 1222
rect 8560 9266 8880 11424
rect 8560 9030 8602 9266
rect 8838 9030 8880 9266
rect 8560 5886 8880 9030
rect 8560 5650 8602 5886
rect 8838 5650 8880 5886
rect 8560 2506 8880 5650
rect 8560 2270 8602 2506
rect 8838 2270 8880 2506
rect 8560 1088 8880 2270
<< via4 >>
rect 2602 8192 2838 8218
rect 2602 8128 2632 8192
rect 2632 8128 2648 8192
rect 2648 8128 2712 8192
rect 2712 8128 2728 8192
rect 2728 8128 2792 8192
rect 2792 8128 2808 8192
rect 2808 8128 2838 8192
rect 2602 7982 2838 8128
rect 2602 4602 2838 4838
rect 2018 3960 2254 4196
rect 1278 2270 1514 2506
rect 2602 1222 2838 1458
rect 3602 9030 3838 9266
rect 3602 5650 3838 5886
rect 3602 2270 3838 2506
rect 5102 9824 5338 9908
rect 5102 9760 5132 9824
rect 5132 9760 5148 9824
rect 5148 9760 5212 9824
rect 5212 9760 5228 9824
rect 5228 9760 5292 9824
rect 5292 9760 5308 9824
rect 5308 9760 5338 9824
rect 5102 9672 5338 9760
rect 5102 6496 5132 6528
rect 5132 6496 5148 6528
rect 5148 6496 5212 6528
rect 5212 6496 5228 6528
rect 5228 6496 5292 6528
rect 5292 6496 5308 6528
rect 5308 6496 5338 6528
rect 5102 6292 5338 6496
rect 5102 2912 5338 3148
rect 6102 10720 6338 10956
rect 6102 7340 6338 7576
rect 6102 3960 6338 4196
rect 7602 8192 7838 8218
rect 7602 8128 7632 8192
rect 7632 8128 7648 8192
rect 7648 8128 7712 8192
rect 7712 8128 7728 8192
rect 7728 8128 7792 8192
rect 7792 8128 7808 8192
rect 7808 8128 7838 8192
rect 7602 7982 7838 8128
rect 7602 4602 7838 4838
rect 7602 1222 7838 1458
rect 8602 9030 8838 9266
rect 8602 5650 8838 5886
rect 8602 2270 8838 2506
<< metal5 >>
rect 920 10956 9844 10998
rect 920 10720 6102 10956
rect 6338 10720 9844 10956
rect 920 10678 9844 10720
rect 920 9908 9844 9950
rect 920 9672 5102 9908
rect 5338 9672 9844 9908
rect 920 9630 9844 9672
rect 920 9266 9844 9308
rect 920 9030 3602 9266
rect 3838 9030 8602 9266
rect 8838 9030 9844 9266
rect 920 8988 9844 9030
rect 920 8218 9844 8260
rect 920 7982 2602 8218
rect 2838 7982 7602 8218
rect 7838 7982 9844 8218
rect 920 7940 9844 7982
rect 920 7576 9844 7618
rect 920 7340 6102 7576
rect 6338 7340 9844 7576
rect 920 7298 9844 7340
rect 920 6528 9844 6570
rect 920 6292 5102 6528
rect 5338 6292 9844 6528
rect 920 6250 9844 6292
rect 920 5886 9844 5928
rect 920 5650 3602 5886
rect 3838 5650 8602 5886
rect 8838 5650 9844 5886
rect 920 5608 9844 5650
rect 920 4838 9844 4880
rect 920 4602 2602 4838
rect 2838 4602 7602 4838
rect 7838 4602 9844 4838
rect 920 4560 9844 4602
rect 920 4196 9844 4238
rect 920 3960 2018 4196
rect 2254 3960 6102 4196
rect 6338 3960 9844 4196
rect 920 3918 9844 3960
rect 920 3148 9844 3190
rect 920 2912 5102 3148
rect 5338 2912 9844 3148
rect 920 2870 9844 2912
rect 920 2506 9844 2548
rect 920 2270 1278 2506
rect 1514 2270 3602 2506
rect 3838 2270 8602 2506
rect 8838 2270 9844 2506
rect 920 2228 9844 2270
rect 920 1458 9844 1500
rect 920 1222 2602 1458
rect 2838 1222 7602 1458
rect 7838 1222 9844 1458
rect 920 1180 9844 1222
use sky130_fd_sc_hd__diode_2  ANTENNA__096__A pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9568 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__098__B
timestamp 1644511149
transform -1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A2
timestamp 1644511149
transform -1 0 8280 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__100__A
timestamp 1644511149
transform -1 0 9568 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A
timestamp 1644511149
transform 1 0 9108 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__102__A
timestamp 1644511149
transform -1 0 8924 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__106__A
timestamp 1644511149
transform 1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A
timestamp 1644511149
transform 1 0 4048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__B
timestamp 1644511149
transform 1 0 2208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__114__A
timestamp 1644511149
transform 1 0 5888 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__B_N
timestamp 1644511149
transform 1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__B
timestamp 1644511149
transform -1 0 3496 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__B_N
timestamp 1644511149
transform -1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__B
timestamp 1644511149
transform 1 0 5244 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__B_N
timestamp 1644511149
transform -1 0 5152 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__B
timestamp 1644511149
transform 1 0 6624 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__B_N
timestamp 1644511149
transform -1 0 7912 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__B
timestamp 1644511149
transform -1 0 4784 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__B_N
timestamp 1644511149
transform 1 0 4140 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__B
timestamp 1644511149
transform -1 0 6348 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__B_N
timestamp 1644511149
transform -1 0 5612 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__B
timestamp 1644511149
transform -1 0 6072 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__B_N
timestamp 1644511149
transform -1 0 1472 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__B
timestamp 1644511149
transform -1 0 9384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__B_N
timestamp 1644511149
transform -1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__B
timestamp 1644511149
transform -1 0 8464 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__B_N
timestamp 1644511149
transform -1 0 3496 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__B
timestamp 1644511149
transform -1 0 8648 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__B_N
timestamp 1644511149
transform -1 0 8096 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__B
timestamp 1644511149
transform -1 0 4600 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__B_N
timestamp 1644511149
transform -1 0 4140 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__172__B
timestamp 1644511149
transform -1 0 4416 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__175__B_N
timestamp 1644511149
transform -1 0 3956 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__177__B
timestamp 1644511149
transform -1 0 3772 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__B_N
timestamp 1644511149
transform -1 0 3588 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__D
timestamp 1644511149
transform -1 0 1564 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__RESET_B
timestamp 1644511149
transform -1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__196__RESET_B
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__RESET_B
timestamp 1644511149
transform -1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__198__RESET_B
timestamp 1644511149
transform -1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__RESET_B
timestamp 1644511149
transform -1 0 1840 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__RESET_B
timestamp 1644511149
transform 1 0 8280 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__RESET_B
timestamp 1644511149
transform 1 0 8464 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__202__RESET_B
timestamp 1644511149
transform 1 0 8648 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__RESET_B
timestamp 1644511149
transform 1 0 8832 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__204__RESET_B
timestamp 1644511149
transform -1 0 8280 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__RESET_B
timestamp 1644511149
transform 1 0 9384 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__RESET_B
timestamp 1644511149
transform -1 0 8464 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__RESET_B
timestamp 1644511149
transform 1 0 9292 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A
timestamp 1644511149
transform -1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A
timestamp 1644511149
transform -1 0 9292 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_clock_A
timestamp 1644511149
transform -1 0 7912 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_serial_load_A
timestamp 1644511149
transform -1 0 8096 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47 pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5244 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_78
timestamp 1644511149
transform 1 0 8096 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_88
timestamp 1644511149
transform 1 0 9016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1644511149
transform 1 0 9476 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_26
timestamp 1644511149
transform 1 0 3312 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_35
timestamp 1644511149
transform 1 0 4140 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_84
timestamp 1644511149
transform 1 0 8648 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_1_93
timestamp 1644511149
transform 1 0 9476 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_47
timestamp 1644511149
transform 1 0 5244 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8556 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_93
timestamp 1644511149
transform 1 0 9476 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_26
timestamp 1644511149
transform 1 0 3312 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_50
timestamp 1644511149
transform 1 0 5520 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_88
timestamp 1644511149
transform 1 0 9016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_26
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp 1644511149
transform 1 0 6348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_26
timestamp 1644511149
transform 1 0 3312 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_85
timestamp 1644511149
transform 1 0 8740 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_3
timestamp 1644511149
transform 1 0 1196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_3
timestamp 1644511149
transform 1 0 1196 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_24
timestamp 1644511149
transform 1 0 3128 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_85
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_3
timestamp 1644511149
transform 1 0 1196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_93
timestamp 1644511149
transform 1 0 9476 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_13_3
timestamp 1644511149
transform 1 0 1196 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_53
timestamp 1644511149
transform 1 0 5796 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1644511149
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 5980 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_3
timestamp 1644511149
transform 1 0 1196 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_32
timestamp 1644511149
transform 1 0 3864 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_93
timestamp 1644511149
transform 1 0 9476 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_79
timestamp 1644511149
transform 1 0 8188 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_3 pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1196 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_7
timestamp 1644511149
transform 1 0 1564 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_13
timestamp 1644511149
transform 1 0 2116 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_42
timestamp 1644511149
transform 1 0 4784 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_46
timestamp 1644511149
transform 1 0 5152 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_18_67
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_0 pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3036 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 9844 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 3036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 9844 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 3036 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 9844 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 3036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 9844 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 3036 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 3036 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 9844 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 3036 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 9844 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 3036 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 9844 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 920 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 9844 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 920 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 9844 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 920 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 9844 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 920 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 9844 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 920 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 9844 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 920 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 9844 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 920 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 9844 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 920 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 9844 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 920 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 9844 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 920 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 9844 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38 pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1644511149
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1644511149
transform 1 0 8188 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1644511149
transform 1 0 5612 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1644511149
transform 1 0 8188 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1644511149
transform 1 0 5612 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1644511149
transform 1 0 8188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1644511149
transform 1 0 5612 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1644511149
transform 1 0 8188 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1644511149
transform 1 0 3496 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1644511149
transform 1 0 6072 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1644511149
transform 1 0 8648 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1644511149
transform 1 0 6072 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1644511149
transform 1 0 3496 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1644511149
transform 1 0 8648 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1644511149
transform 1 0 6072 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1644511149
transform 1 0 3496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1644511149
transform 1 0 8648 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1644511149
transform 1 0 6072 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1644511149
transform 1 0 3496 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1644511149
transform 1 0 8648 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1644511149
transform 1 0 6072 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1644511149
transform 1 0 3496 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1644511149
transform 1 0 8648 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1644511149
transform 1 0 6072 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1644511149
transform 1 0 3496 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1644511149
transform 1 0 6072 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1644511149
transform 1 0 8648 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__or2b_2  _096_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _097_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_2  _098_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_2  _099_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8004 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _100_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8648 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _101_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9292 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _102_
timestamp 1644511149
transform 1 0 8924 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _103_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o31ai_2  _104_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8648 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__o22ai_2  _105_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7360 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _106_
timestamp 1644511149
transform -1 0 9568 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _107_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9568 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  _108_
timestamp 1644511149
transform 1 0 6532 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _109_
timestamp 1644511149
transform -1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _110_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2392 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _111_
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _112_
timestamp 1644511149
transform -1 0 5152 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _113__4
timestamp 1644511149
transform -1 0 2116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _114_
timestamp 1644511149
transform -1 0 5244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _115_
timestamp 1644511149
transform -1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _116_
timestamp 1644511149
transform 1 0 2024 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _117_
timestamp 1644511149
transform -1 0 3864 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _118_
timestamp 1644511149
transform 1 0 2852 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _119_
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _120__5
timestamp 1644511149
transform -1 0 2024 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _121_
timestamp 1644511149
transform 1 0 2668 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _122_
timestamp 1644511149
transform -1 0 3404 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _123_
timestamp 1644511149
transform 1 0 5520 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _124_
timestamp 1644511149
transform 1 0 5428 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _125_
timestamp 1644511149
transform 1 0 5888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _126__6
timestamp 1644511149
transform 1 0 7176 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _127_
timestamp 1644511149
transform 1 0 5152 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _128_
timestamp 1644511149
transform -1 0 7728 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _129_
timestamp 1644511149
transform 1 0 6164 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _130_
timestamp 1644511149
transform 1 0 7912 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _131__7
timestamp 1644511149
transform 1 0 7176 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _132_
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _133_
timestamp 1644511149
transform 1 0 7452 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _134_
timestamp 1644511149
transform 1 0 4508 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _135_
timestamp 1644511149
transform -1 0 6072 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _136__8
timestamp 1644511149
transform 1 0 3864 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _137_
timestamp 1644511149
transform -1 0 4968 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _138_
timestamp 1644511149
transform 1 0 4324 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _139_
timestamp 1644511149
transform 1 0 4968 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _140_
timestamp 1644511149
transform -1 0 6072 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _141_
timestamp 1644511149
transform 1 0 3220 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _142__9
timestamp 1644511149
transform -1 0 6072 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _143_
timestamp 1644511149
transform 1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _144_
timestamp 1644511149
transform -1 0 4232 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _145_
timestamp 1644511149
transform 1 0 1288 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _146_
timestamp 1644511149
transform -1 0 5888 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1644511149
transform 1 0 4232 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _148__10
timestamp 1644511149
transform -1 0 1748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _149_
timestamp 1644511149
transform 1 0 4324 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _150_
timestamp 1644511149
transform -1 0 6440 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _151_
timestamp 1644511149
transform 1 0 7452 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _152_
timestamp 1644511149
transform 1 0 7728 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _153_
timestamp 1644511149
transform -1 0 9568 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _154__11
timestamp 1644511149
transform 1 0 6808 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _155_
timestamp 1644511149
transform 1 0 6164 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _156_
timestamp 1644511149
transform -1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _157_
timestamp 1644511149
transform 1 0 8280 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _158_
timestamp 1644511149
transform -1 0 9016 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _159__12
timestamp 1644511149
transform 1 0 7360 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _160_
timestamp 1644511149
transform 1 0 6808 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _161_
timestamp 1644511149
transform -1 0 9568 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _162_
timestamp 1644511149
transform -1 0 8740 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _163_
timestamp 1644511149
transform 1 0 7636 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _164__13
timestamp 1644511149
transform -1 0 5060 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _165_
timestamp 1644511149
transform 1 0 7084 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _166_
timestamp 1644511149
transform -1 0 8188 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _167_
timestamp 1644511149
transform 1 0 5060 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _168_
timestamp 1644511149
transform 1 0 4508 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _169__1
timestamp 1644511149
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _170_
timestamp 1644511149
transform -1 0 4784 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _171_
timestamp 1644511149
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _172_
timestamp 1644511149
transform 1 0 5704 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _173_
timestamp 1644511149
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _174__2
timestamp 1644511149
transform -1 0 3772 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _175_
timestamp 1644511149
transform -1 0 5428 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _176_
timestamp 1644511149
transform 1 0 3404 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _177_
timestamp 1644511149
transform 1 0 3956 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _178_
timestamp 1644511149
transform -1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _179__3
timestamp 1644511149
transform 1 0 5336 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _180_
timestamp 1644511149
transform 1 0 5704 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  _181_
timestamp 1644511149
transform 1 0 5336 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__dfbbn_2  _182_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1748 0 -1 10880
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _183_
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _184_
timestamp 1644511149
transform -1 0 8372 0 1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _185_
timestamp 1644511149
transform 1 0 6808 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _186_
timestamp 1644511149
transform 1 0 3404 0 -1 9792
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _187_
timestamp 1644511149
transform 1 0 3220 0 -1 6528
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _188_
timestamp 1644511149
transform 1 0 3496 0 -1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _189_
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _190_
timestamp 1644511149
transform 1 0 6440 0 1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _191_
timestamp 1644511149
transform 1 0 6348 0 1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _192_
timestamp 1644511149
transform 1 0 3680 0 -1 3264
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _193_
timestamp 1644511149
transform 1 0 4416 0 -1 4352
box -38 -48 2614 592
use sky130_fd_sc_hd__dfbbn_2  _194_
timestamp 1644511149
transform 1 0 5980 0 1 2176
box -38 -48 2614 592
use sky130_fd_sc_hd__dfrtp_2  _195_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 1196 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _196_
timestamp 1644511149
transform -1 0 3496 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _197_
timestamp 1644511149
transform -1 0 3128 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _198_
timestamp 1644511149
transform 1 0 1288 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _199_
timestamp 1644511149
transform 1 0 1564 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _200_
timestamp 1644511149
transform 1 0 3312 0 1 1088
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _201_
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _202_
timestamp 1644511149
transform 1 0 4600 0 -1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _203_
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _204_
timestamp 1644511149
transform -1 0 8096 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _205_
timestamp 1644511149
transform -1 0 9200 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _206_
timestamp 1644511149
transform 1 0 6072 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _207_
timestamp 1644511149
transform 1 0 7360 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_2  _208_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9200 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _209_
timestamp 1644511149
transform 1 0 8280 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _210_
timestamp 1644511149
transform 1 0 8280 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__ebufn_2  _211_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9476 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__049_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4232 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__077_
timestamp 1644511149
transform -1 0 5796 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock
timestamp 1644511149
transform -1 0 7084 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_load
timestamp 1644511149
transform -1 0 7912 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__049_ pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6992 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0__077_
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_clock
timestamp 1644511149
transform -1 0 3956 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_serial_load
timestamp 1644511149
transform -1 0 5244 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__049_
timestamp 1644511149
transform -1 0 4232 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0__077_
timestamp 1644511149
transform 1 0 6808 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_clock
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_serial_load
timestamp 1644511149
transform -1 0 6532 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  const_source pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9476 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6532 0 -1 2176
box -38 -48 1694 592
use gpio_logic_high  gpio_logic_high
timestamp 0
transform 1 0 1196 0 1 1680
box -38 -48 1418 2768
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold1 pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold2
timestamp 1644511149
transform 1 0 3404 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold3
timestamp 1644511149
transform -1 0 2024 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold4
timestamp 1644511149
transform -1 0 2024 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold5
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold6
timestamp 1644511149
transform -1 0 4324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold7 pdks_with_sram/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9016 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold8
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold9
timestamp 1644511149
transform -1 0 8648 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold10
timestamp 1644511149
transform -1 0 9568 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold11
timestamp 1644511149
transform 1 0 4324 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold12
timestamp 1644511149
transform 1 0 5060 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold13
timestamp 1644511149
transform 1 0 4140 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold14
timestamp 1644511149
transform -1 0 4140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold15
timestamp 1644511149
transform 1 0 2024 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold16
timestamp 1644511149
transform 1 0 2760 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold17
timestamp 1644511149
transform 1 0 2024 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold18
timestamp 1644511149
transform -1 0 3496 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold19
timestamp 1644511149
transform 1 0 4324 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold20
timestamp 1644511149
transform 1 0 5060 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold21
timestamp 1644511149
transform -1 0 9476 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold22
timestamp 1644511149
transform 1 0 6532 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold23
timestamp 1644511149
transform -1 0 9384 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold24
timestamp 1644511149
transform -1 0 7176 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold25
timestamp 1644511149
transform 1 0 5704 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__clkdlybuf4s25_1  hold26
timestamp 1644511149
transform 1 0 7176 0 1 1088
box -38 -48 774 592
<< labels >>
rlabel metal2 s 938 12200 994 13000 6 gpio_defaults[0]
port 0 nsew signal input
rlabel metal2 s 5538 12200 5594 13000 6 gpio_defaults[10]
port 1 nsew signal input
rlabel metal2 s 5998 12200 6054 13000 6 gpio_defaults[11]
port 2 nsew signal input
rlabel metal2 s 6458 12200 6514 13000 6 gpio_defaults[12]
port 3 nsew signal input
rlabel metal2 s 1398 12200 1454 13000 6 gpio_defaults[1]
port 4 nsew signal input
rlabel metal2 s 1858 12200 1914 13000 6 gpio_defaults[2]
port 5 nsew signal input
rlabel metal2 s 2318 12200 2374 13000 6 gpio_defaults[3]
port 6 nsew signal input
rlabel metal2 s 2778 12200 2834 13000 6 gpio_defaults[4]
port 7 nsew signal input
rlabel metal2 s 3238 12200 3294 13000 6 gpio_defaults[5]
port 8 nsew signal input
rlabel metal2 s 3698 12200 3754 13000 6 gpio_defaults[6]
port 9 nsew signal input
rlabel metal2 s 4158 12200 4214 13000 6 gpio_defaults[7]
port 10 nsew signal input
rlabel metal2 s 4618 12200 4674 13000 6 gpio_defaults[8]
port 11 nsew signal input
rlabel metal2 s 5078 12200 5134 13000 6 gpio_defaults[9]
port 12 nsew signal input
rlabel metal3 s 14000 824 34000 944 6 mgmt_gpio_in
port 13 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 14 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 15 nsew signal input
rlabel metal3 s 14000 1232 34000 1352 6 one
port 16 nsew signal tristate
rlabel metal3 s 14000 2456 34000 2576 6 pad_gpio_ana_en
port 17 nsew signal tristate
rlabel metal3 s 14000 2864 34000 2984 6 pad_gpio_ana_pol
port 18 nsew signal tristate
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_sel
port 19 nsew signal tristate
rlabel metal3 s 14000 3680 34000 3800 6 pad_gpio_dm[0]
port 20 nsew signal tristate
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[1]
port 21 nsew signal tristate
rlabel metal3 s 14000 4496 34000 4616 6 pad_gpio_dm[2]
port 22 nsew signal tristate
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_holdover
port 23 nsew signal tristate
rlabel metal3 s 14000 5312 34000 5432 6 pad_gpio_ib_mode_sel
port 24 nsew signal tristate
rlabel metal3 s 14000 5720 34000 5840 6 pad_gpio_in
port 25 nsew signal input
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_inenb
port 26 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_out
port 27 nsew signal tristate
rlabel metal3 s 14000 6944 34000 7064 6 pad_gpio_outenb
port 28 nsew signal tristate
rlabel metal3 s 14000 7352 34000 7472 6 pad_gpio_slow_sel
port 29 nsew signal tristate
rlabel metal3 s 14000 7760 34000 7880 6 pad_gpio_vtrip_sel
port 30 nsew signal tristate
rlabel metal3 s 14000 8168 34000 8288 6 resetn
port 31 nsew signal input
rlabel metal3 s 14000 8576 34000 8696 6 resetn_out
port 32 nsew signal tristate
rlabel metal3 s 14000 8984 34000 9104 6 serial_clock
port 33 nsew signal input
rlabel metal3 s 14000 9392 34000 9512 6 serial_clock_out
port 34 nsew signal tristate
rlabel metal3 s 14000 9800 34000 9920 6 serial_data_in
port 35 nsew signal input
rlabel metal3 s 14000 10208 34000 10328 6 serial_data_out
port 36 nsew signal tristate
rlabel metal3 s 14000 10616 34000 10736 6 serial_load
port 37 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_load_out
port 38 nsew signal tristate
rlabel metal3 s 14000 11432 34000 11552 6 user_gpio_in
port 39 nsew signal tristate
rlabel metal3 s 14000 11840 34000 11960 6 user_gpio_oeb
port 40 nsew signal input
rlabel metal3 s 14000 12248 34000 12368 6 user_gpio_out
port 41 nsew signal input
rlabel metal5 s 920 1180 9844 1500 6 vccd
port 42 nsew power input
rlabel metal5 s 920 4560 9844 4880 6 vccd
port 42 nsew power input
rlabel metal5 s 920 7940 9844 8260 6 vccd
port 42 nsew power input
rlabel metal4 s 2560 1088 2880 11472 6 vccd
port 42 nsew power input
rlabel metal4 s 7560 1040 7880 11472 6 vccd
port 42 nsew power input
rlabel metal5 s 920 2228 9844 2548 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 5608 9844 5928 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 8988 9844 9308 6 vccd1
port 43 nsew power input
rlabel metal4 s 3560 1088 3880 11424 6 vccd1
port 43 nsew power input
rlabel metal4 s 8560 1088 8880 11424 6 vccd1
port 43 nsew power input
rlabel metal5 s 920 2870 9844 3190 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 6250 9844 6570 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 9630 9844 9950 6 vssd
port 44 nsew ground input
rlabel metal4 s 5060 1040 5380 11472 6 vssd
port 44 nsew ground input
rlabel metal5 s 920 3918 9844 4238 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 7298 9844 7618 6 vssd1
port 45 nsew ground input
rlabel metal5 s 920 10678 9844 10998 6 vssd1
port 45 nsew ground input
rlabel metal4 s 6060 1088 6380 11424 6 vssd1
port 45 nsew ground input
rlabel metal3 s 14000 416 34000 536 6 zero
port 46 nsew signal tristate
<< properties >>
string FIXED_BBOX 0 0 34000 13000
<< end >>
